magic
tech sky130A
magscale 1 2
timestamp 1716907293
<< nwell >>
rect -496 -519 496 519
<< pmoslvt >>
rect -300 -300 300 300
<< pdiff >>
rect -358 288 -300 300
rect -358 -288 -346 288
rect -312 -288 -300 288
rect -358 -300 -300 -288
rect 300 288 358 300
rect 300 -288 312 288
rect 346 -288 358 288
rect 300 -300 358 -288
<< pdiffc >>
rect -346 -288 -312 288
rect 312 -288 346 288
<< nsubdiff >>
rect -460 449 -364 483
rect 364 449 460 483
rect -460 387 -426 449
rect 426 387 460 449
rect -460 -449 -426 -387
rect 426 -449 460 -387
rect -460 -483 -364 -449
rect 364 -483 460 -449
<< nsubdiffcont >>
rect -364 449 364 483
rect -460 -387 -426 387
rect 426 -387 460 387
rect -364 -483 364 -449
<< poly >>
rect -300 381 300 397
rect -300 347 -284 381
rect 284 347 300 381
rect -300 300 300 347
rect -300 -347 300 -300
rect -300 -381 -284 -347
rect 284 -381 300 -347
rect -300 -397 300 -381
<< polycont >>
rect -284 347 284 381
rect -284 -381 284 -347
<< locali >>
rect -460 449 -364 483
rect 364 449 460 483
rect -460 387 -426 449
rect 426 387 460 449
rect -300 347 -284 381
rect 284 347 300 381
rect -346 288 -312 304
rect -346 -304 -312 -288
rect 312 288 346 304
rect 312 -304 346 -288
rect -300 -381 -284 -347
rect 284 -381 300 -347
rect -460 -449 -426 -387
rect 426 -449 460 -387
rect -460 -483 -364 -449
rect 364 -483 460 -449
<< viali >>
rect -284 347 284 381
rect -346 -288 -312 288
rect 312 -288 346 288
rect -284 -381 284 -347
<< metal1 >>
rect -296 381 296 387
rect -296 347 -284 381
rect 284 347 296 381
rect -296 341 296 347
rect -352 288 -306 300
rect -352 -288 -346 288
rect -312 -288 -306 288
rect -352 -300 -306 -288
rect 306 288 352 300
rect 306 -288 312 288
rect 346 -288 352 288
rect 306 -300 352 -288
rect -296 -347 296 -341
rect -296 -381 -284 -347
rect 284 -381 296 -347
rect -296 -387 296 -381
<< properties >>
string FIXED_BBOX -443 -466 443 466
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 3.0 l 3.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

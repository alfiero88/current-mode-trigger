magic
tech sky130A
magscale 1 2
timestamp 1716907293
<< error_p >>
rect -351 381 -289 387
rect -223 381 -161 387
rect -95 381 -33 387
rect 33 381 95 387
rect 161 381 223 387
rect 289 381 351 387
rect -351 347 -339 381
rect -223 347 -211 381
rect -95 347 -83 381
rect 33 347 45 381
rect 161 347 173 381
rect 289 347 301 381
rect -351 341 -289 347
rect -223 341 -161 347
rect -95 341 -33 347
rect 33 341 95 347
rect 161 341 223 347
rect 289 341 351 347
rect -351 -347 -289 -341
rect -223 -347 -161 -341
rect -95 -347 -33 -341
rect 33 -347 95 -341
rect 161 -347 223 -341
rect 289 -347 351 -341
rect -351 -381 -339 -347
rect -223 -381 -211 -347
rect -95 -381 -83 -347
rect 33 -381 45 -347
rect 161 -381 173 -347
rect 289 -381 301 -347
rect -351 -387 -289 -381
rect -223 -387 -161 -381
rect -95 -387 -33 -381
rect 33 -387 95 -381
rect 161 -387 223 -381
rect 289 -387 351 -381
<< nwell >>
rect -551 -519 551 519
<< pmoslvt >>
rect -355 -300 -285 300
rect -227 -300 -157 300
rect -99 -300 -29 300
rect 29 -300 99 300
rect 157 -300 227 300
rect 285 -300 355 300
<< pdiff >>
rect -413 288 -355 300
rect -413 -288 -401 288
rect -367 -288 -355 288
rect -413 -300 -355 -288
rect -285 288 -227 300
rect -285 -288 -273 288
rect -239 -288 -227 288
rect -285 -300 -227 -288
rect -157 288 -99 300
rect -157 -288 -145 288
rect -111 -288 -99 288
rect -157 -300 -99 -288
rect -29 288 29 300
rect -29 -288 -17 288
rect 17 -288 29 288
rect -29 -300 29 -288
rect 99 288 157 300
rect 99 -288 111 288
rect 145 -288 157 288
rect 99 -300 157 -288
rect 227 288 285 300
rect 227 -288 239 288
rect 273 -288 285 288
rect 227 -300 285 -288
rect 355 288 413 300
rect 355 -288 367 288
rect 401 -288 413 288
rect 355 -300 413 -288
<< pdiffc >>
rect -401 -288 -367 288
rect -273 -288 -239 288
rect -145 -288 -111 288
rect -17 -288 17 288
rect 111 -288 145 288
rect 239 -288 273 288
rect 367 -288 401 288
<< nsubdiff >>
rect -515 449 -419 483
rect 419 449 515 483
rect -515 387 -481 449
rect 481 387 515 449
rect -515 -449 -481 -387
rect 481 -449 515 -387
rect -515 -483 -419 -449
rect 419 -483 515 -449
<< nsubdiffcont >>
rect -419 449 419 483
rect -515 -387 -481 387
rect 481 -387 515 387
rect -419 -483 419 -449
<< poly >>
rect -355 381 -285 397
rect -355 347 -339 381
rect -301 347 -285 381
rect -355 300 -285 347
rect -227 381 -157 397
rect -227 347 -211 381
rect -173 347 -157 381
rect -227 300 -157 347
rect -99 381 -29 397
rect -99 347 -83 381
rect -45 347 -29 381
rect -99 300 -29 347
rect 29 381 99 397
rect 29 347 45 381
rect 83 347 99 381
rect 29 300 99 347
rect 157 381 227 397
rect 157 347 173 381
rect 211 347 227 381
rect 157 300 227 347
rect 285 381 355 397
rect 285 347 301 381
rect 339 347 355 381
rect 285 300 355 347
rect -355 -347 -285 -300
rect -355 -381 -339 -347
rect -301 -381 -285 -347
rect -355 -397 -285 -381
rect -227 -347 -157 -300
rect -227 -381 -211 -347
rect -173 -381 -157 -347
rect -227 -397 -157 -381
rect -99 -347 -29 -300
rect -99 -381 -83 -347
rect -45 -381 -29 -347
rect -99 -397 -29 -381
rect 29 -347 99 -300
rect 29 -381 45 -347
rect 83 -381 99 -347
rect 29 -397 99 -381
rect 157 -347 227 -300
rect 157 -381 173 -347
rect 211 -381 227 -347
rect 157 -397 227 -381
rect 285 -347 355 -300
rect 285 -381 301 -347
rect 339 -381 355 -347
rect 285 -397 355 -381
<< polycont >>
rect -339 347 -301 381
rect -211 347 -173 381
rect -83 347 -45 381
rect 45 347 83 381
rect 173 347 211 381
rect 301 347 339 381
rect -339 -381 -301 -347
rect -211 -381 -173 -347
rect -83 -381 -45 -347
rect 45 -381 83 -347
rect 173 -381 211 -347
rect 301 -381 339 -347
<< locali >>
rect -515 449 -419 483
rect 419 449 515 483
rect -515 387 -481 449
rect 481 387 515 449
rect -355 347 -339 381
rect -301 347 -285 381
rect -227 347 -211 381
rect -173 347 -157 381
rect -99 347 -83 381
rect -45 347 -29 381
rect 29 347 45 381
rect 83 347 99 381
rect 157 347 173 381
rect 211 347 227 381
rect 285 347 301 381
rect 339 347 355 381
rect -401 288 -367 304
rect -401 -304 -367 -288
rect -273 288 -239 304
rect -273 -304 -239 -288
rect -145 288 -111 304
rect -145 -304 -111 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 111 288 145 304
rect 111 -304 145 -288
rect 239 288 273 304
rect 239 -304 273 -288
rect 367 288 401 304
rect 367 -304 401 -288
rect -355 -381 -339 -347
rect -301 -381 -285 -347
rect -227 -381 -211 -347
rect -173 -381 -157 -347
rect -99 -381 -83 -347
rect -45 -381 -29 -347
rect 29 -381 45 -347
rect 83 -381 99 -347
rect 157 -381 173 -347
rect 211 -381 227 -347
rect 285 -381 301 -347
rect 339 -381 355 -347
rect -515 -449 -481 -387
rect 481 -449 515 -387
rect -515 -483 -419 -449
rect 419 -483 515 -449
<< viali >>
rect -339 347 -301 381
rect -211 347 -173 381
rect -83 347 -45 381
rect 45 347 83 381
rect 173 347 211 381
rect 301 347 339 381
rect -401 -288 -367 288
rect -273 -288 -239 288
rect -145 -288 -111 288
rect -17 -288 17 288
rect 111 -288 145 288
rect 239 -288 273 288
rect 367 -288 401 288
rect -339 -381 -301 -347
rect -211 -381 -173 -347
rect -83 -381 -45 -347
rect 45 -381 83 -347
rect 173 -381 211 -347
rect 301 -381 339 -347
<< metal1 >>
rect -351 381 -289 387
rect -351 347 -339 381
rect -301 347 -289 381
rect -351 341 -289 347
rect -223 381 -161 387
rect -223 347 -211 381
rect -173 347 -161 381
rect -223 341 -161 347
rect -95 381 -33 387
rect -95 347 -83 381
rect -45 347 -33 381
rect -95 341 -33 347
rect 33 381 95 387
rect 33 347 45 381
rect 83 347 95 381
rect 33 341 95 347
rect 161 381 223 387
rect 161 347 173 381
rect 211 347 223 381
rect 161 341 223 347
rect 289 381 351 387
rect 289 347 301 381
rect 339 347 351 381
rect 289 341 351 347
rect -407 288 -361 300
rect -407 -288 -401 288
rect -367 -288 -361 288
rect -407 -300 -361 -288
rect -279 288 -233 300
rect -279 -288 -273 288
rect -239 -288 -233 288
rect -279 -300 -233 -288
rect -151 288 -105 300
rect -151 -288 -145 288
rect -111 -288 -105 288
rect -151 -300 -105 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 105 288 151 300
rect 105 -288 111 288
rect 145 -288 151 288
rect 105 -300 151 -288
rect 233 288 279 300
rect 233 -288 239 288
rect 273 -288 279 288
rect 233 -300 279 -288
rect 361 288 407 300
rect 361 -288 367 288
rect 401 -288 407 288
rect 361 -300 407 -288
rect -351 -347 -289 -341
rect -351 -381 -339 -347
rect -301 -381 -289 -347
rect -351 -387 -289 -381
rect -223 -347 -161 -341
rect -223 -381 -211 -347
rect -173 -381 -161 -347
rect -223 -387 -161 -381
rect -95 -347 -33 -341
rect -95 -381 -83 -347
rect -45 -381 -33 -347
rect -95 -387 -33 -381
rect 33 -347 95 -341
rect 33 -381 45 -347
rect 83 -381 95 -347
rect 33 -387 95 -381
rect 161 -347 223 -341
rect 161 -381 173 -347
rect 211 -381 223 -347
rect 161 -387 223 -381
rect 289 -347 351 -341
rect 289 -381 301 -347
rect 339 -381 351 -347
rect 289 -387 351 -381
<< properties >>
string FIXED_BBOX -498 -466 498 466
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 3.0 l 0.35 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

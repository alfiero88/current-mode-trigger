magic
tech sky130A
magscale 1 2
timestamp 1716907293
<< error_p >>
rect -159 281 -97 287
rect -31 281 31 287
rect 97 281 159 287
rect -159 247 -147 281
rect -31 247 -19 281
rect 97 247 109 281
rect -159 241 -97 247
rect -31 241 31 247
rect 97 241 159 247
rect -159 -247 -97 -241
rect -31 -247 31 -241
rect 97 -247 159 -241
rect -159 -281 -147 -247
rect -31 -281 -19 -247
rect 97 -281 109 -247
rect -159 -287 -97 -281
rect -31 -287 31 -281
rect 97 -287 159 -281
<< nwell >>
rect -359 -419 359 419
<< pmoslvt >>
rect -163 -200 -93 200
rect -35 -200 35 200
rect 93 -200 163 200
<< pdiff >>
rect -221 188 -163 200
rect -221 -188 -209 188
rect -175 -188 -163 188
rect -221 -200 -163 -188
rect -93 188 -35 200
rect -93 -188 -81 188
rect -47 -188 -35 188
rect -93 -200 -35 -188
rect 35 188 93 200
rect 35 -188 47 188
rect 81 -188 93 188
rect 35 -200 93 -188
rect 163 188 221 200
rect 163 -188 175 188
rect 209 -188 221 188
rect 163 -200 221 -188
<< pdiffc >>
rect -209 -188 -175 188
rect -81 -188 -47 188
rect 47 -188 81 188
rect 175 -188 209 188
<< nsubdiff >>
rect -323 349 -227 383
rect 227 349 323 383
rect -323 287 -289 349
rect 289 287 323 349
rect -323 -349 -289 -287
rect 289 -349 323 -287
rect -323 -383 -227 -349
rect 227 -383 323 -349
<< nsubdiffcont >>
rect -227 349 227 383
rect -323 -287 -289 287
rect 289 -287 323 287
rect -227 -383 227 -349
<< poly >>
rect -163 281 -93 297
rect -163 247 -147 281
rect -109 247 -93 281
rect -163 200 -93 247
rect -35 281 35 297
rect -35 247 -19 281
rect 19 247 35 281
rect -35 200 35 247
rect 93 281 163 297
rect 93 247 109 281
rect 147 247 163 281
rect 93 200 163 247
rect -163 -247 -93 -200
rect -163 -281 -147 -247
rect -109 -281 -93 -247
rect -163 -297 -93 -281
rect -35 -247 35 -200
rect -35 -281 -19 -247
rect 19 -281 35 -247
rect -35 -297 35 -281
rect 93 -247 163 -200
rect 93 -281 109 -247
rect 147 -281 163 -247
rect 93 -297 163 -281
<< polycont >>
rect -147 247 -109 281
rect -19 247 19 281
rect 109 247 147 281
rect -147 -281 -109 -247
rect -19 -281 19 -247
rect 109 -281 147 -247
<< locali >>
rect -323 349 -227 383
rect 227 349 323 383
rect -323 287 -289 349
rect 289 287 323 349
rect -163 247 -147 281
rect -109 247 -93 281
rect -35 247 -19 281
rect 19 247 35 281
rect 93 247 109 281
rect 147 247 163 281
rect -209 188 -175 204
rect -209 -204 -175 -188
rect -81 188 -47 204
rect -81 -204 -47 -188
rect 47 188 81 204
rect 47 -204 81 -188
rect 175 188 209 204
rect 175 -204 209 -188
rect -163 -281 -147 -247
rect -109 -281 -93 -247
rect -35 -281 -19 -247
rect 19 -281 35 -247
rect 93 -281 109 -247
rect 147 -281 163 -247
rect -323 -349 -289 -287
rect 289 -349 323 -287
rect -323 -383 -227 -349
rect 227 -383 323 -349
<< viali >>
rect -147 247 -109 281
rect -19 247 19 281
rect 109 247 147 281
rect -209 -188 -175 188
rect -81 -188 -47 188
rect 47 -188 81 188
rect 175 -188 209 188
rect -147 -281 -109 -247
rect -19 -281 19 -247
rect 109 -281 147 -247
<< metal1 >>
rect -159 281 -97 287
rect -159 247 -147 281
rect -109 247 -97 281
rect -159 241 -97 247
rect -31 281 31 287
rect -31 247 -19 281
rect 19 247 31 281
rect -31 241 31 247
rect 97 281 159 287
rect 97 247 109 281
rect 147 247 159 281
rect 97 241 159 247
rect -215 188 -169 200
rect -215 -188 -209 188
rect -175 -188 -169 188
rect -215 -200 -169 -188
rect -87 188 -41 200
rect -87 -188 -81 188
rect -47 -188 -41 188
rect -87 -200 -41 -188
rect 41 188 87 200
rect 41 -188 47 188
rect 81 -188 87 188
rect 41 -200 87 -188
rect 169 188 215 200
rect 169 -188 175 188
rect 209 -188 215 188
rect 169 -200 215 -188
rect -159 -247 -97 -241
rect -159 -281 -147 -247
rect -109 -281 -97 -247
rect -159 -287 -97 -281
rect -31 -247 31 -241
rect -31 -281 -19 -247
rect 19 -281 31 -247
rect -31 -287 31 -281
rect 97 -247 159 -241
rect 97 -281 109 -247
rect 147 -281 159 -247
rect 97 -287 159 -281
<< properties >>
string FIXED_BBOX -306 -366 306 366
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 2.0 l 0.35 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1716907293
<< nwell >>
rect -3128 -419 3128 419
<< pmoslvt >>
rect -2932 -200 -2332 200
rect -2274 -200 -1674 200
rect -1616 -200 -1016 200
rect -958 -200 -358 200
rect -300 -200 300 200
rect 358 -200 958 200
rect 1016 -200 1616 200
rect 1674 -200 2274 200
rect 2332 -200 2932 200
<< pdiff >>
rect -2990 188 -2932 200
rect -2990 -188 -2978 188
rect -2944 -188 -2932 188
rect -2990 -200 -2932 -188
rect -2332 188 -2274 200
rect -2332 -188 -2320 188
rect -2286 -188 -2274 188
rect -2332 -200 -2274 -188
rect -1674 188 -1616 200
rect -1674 -188 -1662 188
rect -1628 -188 -1616 188
rect -1674 -200 -1616 -188
rect -1016 188 -958 200
rect -1016 -188 -1004 188
rect -970 -188 -958 188
rect -1016 -200 -958 -188
rect -358 188 -300 200
rect -358 -188 -346 188
rect -312 -188 -300 188
rect -358 -200 -300 -188
rect 300 188 358 200
rect 300 -188 312 188
rect 346 -188 358 188
rect 300 -200 358 -188
rect 958 188 1016 200
rect 958 -188 970 188
rect 1004 -188 1016 188
rect 958 -200 1016 -188
rect 1616 188 1674 200
rect 1616 -188 1628 188
rect 1662 -188 1674 188
rect 1616 -200 1674 -188
rect 2274 188 2332 200
rect 2274 -188 2286 188
rect 2320 -188 2332 188
rect 2274 -200 2332 -188
rect 2932 188 2990 200
rect 2932 -188 2944 188
rect 2978 -188 2990 188
rect 2932 -200 2990 -188
<< pdiffc >>
rect -2978 -188 -2944 188
rect -2320 -188 -2286 188
rect -1662 -188 -1628 188
rect -1004 -188 -970 188
rect -346 -188 -312 188
rect 312 -188 346 188
rect 970 -188 1004 188
rect 1628 -188 1662 188
rect 2286 -188 2320 188
rect 2944 -188 2978 188
<< nsubdiff >>
rect -3092 349 -2996 383
rect 2996 349 3092 383
rect -3092 287 -3058 349
rect 3058 287 3092 349
rect -3092 -349 -3058 -287
rect 3058 -349 3092 -287
rect -3092 -383 -2996 -349
rect 2996 -383 3092 -349
<< nsubdiffcont >>
rect -2996 349 2996 383
rect -3092 -287 -3058 287
rect 3058 -287 3092 287
rect -2996 -383 2996 -349
<< poly >>
rect -2932 281 -2332 297
rect -2932 247 -2916 281
rect -2348 247 -2332 281
rect -2932 200 -2332 247
rect -2274 281 -1674 297
rect -2274 247 -2258 281
rect -1690 247 -1674 281
rect -2274 200 -1674 247
rect -1616 281 -1016 297
rect -1616 247 -1600 281
rect -1032 247 -1016 281
rect -1616 200 -1016 247
rect -958 281 -358 297
rect -958 247 -942 281
rect -374 247 -358 281
rect -958 200 -358 247
rect -300 281 300 297
rect -300 247 -284 281
rect 284 247 300 281
rect -300 200 300 247
rect 358 281 958 297
rect 358 247 374 281
rect 942 247 958 281
rect 358 200 958 247
rect 1016 281 1616 297
rect 1016 247 1032 281
rect 1600 247 1616 281
rect 1016 200 1616 247
rect 1674 281 2274 297
rect 1674 247 1690 281
rect 2258 247 2274 281
rect 1674 200 2274 247
rect 2332 281 2932 297
rect 2332 247 2348 281
rect 2916 247 2932 281
rect 2332 200 2932 247
rect -2932 -247 -2332 -200
rect -2932 -281 -2916 -247
rect -2348 -281 -2332 -247
rect -2932 -297 -2332 -281
rect -2274 -247 -1674 -200
rect -2274 -281 -2258 -247
rect -1690 -281 -1674 -247
rect -2274 -297 -1674 -281
rect -1616 -247 -1016 -200
rect -1616 -281 -1600 -247
rect -1032 -281 -1016 -247
rect -1616 -297 -1016 -281
rect -958 -247 -358 -200
rect -958 -281 -942 -247
rect -374 -281 -358 -247
rect -958 -297 -358 -281
rect -300 -247 300 -200
rect -300 -281 -284 -247
rect 284 -281 300 -247
rect -300 -297 300 -281
rect 358 -247 958 -200
rect 358 -281 374 -247
rect 942 -281 958 -247
rect 358 -297 958 -281
rect 1016 -247 1616 -200
rect 1016 -281 1032 -247
rect 1600 -281 1616 -247
rect 1016 -297 1616 -281
rect 1674 -247 2274 -200
rect 1674 -281 1690 -247
rect 2258 -281 2274 -247
rect 1674 -297 2274 -281
rect 2332 -247 2932 -200
rect 2332 -281 2348 -247
rect 2916 -281 2932 -247
rect 2332 -297 2932 -281
<< polycont >>
rect -2916 247 -2348 281
rect -2258 247 -1690 281
rect -1600 247 -1032 281
rect -942 247 -374 281
rect -284 247 284 281
rect 374 247 942 281
rect 1032 247 1600 281
rect 1690 247 2258 281
rect 2348 247 2916 281
rect -2916 -281 -2348 -247
rect -2258 -281 -1690 -247
rect -1600 -281 -1032 -247
rect -942 -281 -374 -247
rect -284 -281 284 -247
rect 374 -281 942 -247
rect 1032 -281 1600 -247
rect 1690 -281 2258 -247
rect 2348 -281 2916 -247
<< locali >>
rect -3092 349 -2996 383
rect 2996 349 3092 383
rect -3092 287 -3058 349
rect 3058 287 3092 349
rect -2932 247 -2916 281
rect -2348 247 -2332 281
rect -2274 247 -2258 281
rect -1690 247 -1674 281
rect -1616 247 -1600 281
rect -1032 247 -1016 281
rect -958 247 -942 281
rect -374 247 -358 281
rect -300 247 -284 281
rect 284 247 300 281
rect 358 247 374 281
rect 942 247 958 281
rect 1016 247 1032 281
rect 1600 247 1616 281
rect 1674 247 1690 281
rect 2258 247 2274 281
rect 2332 247 2348 281
rect 2916 247 2932 281
rect -2978 188 -2944 204
rect -2978 -204 -2944 -188
rect -2320 188 -2286 204
rect -2320 -204 -2286 -188
rect -1662 188 -1628 204
rect -1662 -204 -1628 -188
rect -1004 188 -970 204
rect -1004 -204 -970 -188
rect -346 188 -312 204
rect -346 -204 -312 -188
rect 312 188 346 204
rect 312 -204 346 -188
rect 970 188 1004 204
rect 970 -204 1004 -188
rect 1628 188 1662 204
rect 1628 -204 1662 -188
rect 2286 188 2320 204
rect 2286 -204 2320 -188
rect 2944 188 2978 204
rect 2944 -204 2978 -188
rect -2932 -281 -2916 -247
rect -2348 -281 -2332 -247
rect -2274 -281 -2258 -247
rect -1690 -281 -1674 -247
rect -1616 -281 -1600 -247
rect -1032 -281 -1016 -247
rect -958 -281 -942 -247
rect -374 -281 -358 -247
rect -300 -281 -284 -247
rect 284 -281 300 -247
rect 358 -281 374 -247
rect 942 -281 958 -247
rect 1016 -281 1032 -247
rect 1600 -281 1616 -247
rect 1674 -281 1690 -247
rect 2258 -281 2274 -247
rect 2332 -281 2348 -247
rect 2916 -281 2932 -247
rect -3092 -349 -3058 -287
rect 3058 -349 3092 -287
rect -3092 -383 -2996 -349
rect 2996 -383 3092 -349
<< viali >>
rect -2916 247 -2348 281
rect -2258 247 -1690 281
rect -1600 247 -1032 281
rect -942 247 -374 281
rect -284 247 284 281
rect 374 247 942 281
rect 1032 247 1600 281
rect 1690 247 2258 281
rect 2348 247 2916 281
rect -2978 -188 -2944 188
rect -2320 -188 -2286 188
rect -1662 -188 -1628 188
rect -1004 -188 -970 188
rect -346 -188 -312 188
rect 312 -188 346 188
rect 970 -188 1004 188
rect 1628 -188 1662 188
rect 2286 -188 2320 188
rect 2944 -188 2978 188
rect -2916 -281 -2348 -247
rect -2258 -281 -1690 -247
rect -1600 -281 -1032 -247
rect -942 -281 -374 -247
rect -284 -281 284 -247
rect 374 -281 942 -247
rect 1032 -281 1600 -247
rect 1690 -281 2258 -247
rect 2348 -281 2916 -247
<< metal1 >>
rect -2928 281 -2336 287
rect -2928 247 -2916 281
rect -2348 247 -2336 281
rect -2928 241 -2336 247
rect -2270 281 -1678 287
rect -2270 247 -2258 281
rect -1690 247 -1678 281
rect -2270 241 -1678 247
rect -1612 281 -1020 287
rect -1612 247 -1600 281
rect -1032 247 -1020 281
rect -1612 241 -1020 247
rect -954 281 -362 287
rect -954 247 -942 281
rect -374 247 -362 281
rect -954 241 -362 247
rect -296 281 296 287
rect -296 247 -284 281
rect 284 247 296 281
rect -296 241 296 247
rect 362 281 954 287
rect 362 247 374 281
rect 942 247 954 281
rect 362 241 954 247
rect 1020 281 1612 287
rect 1020 247 1032 281
rect 1600 247 1612 281
rect 1020 241 1612 247
rect 1678 281 2270 287
rect 1678 247 1690 281
rect 2258 247 2270 281
rect 1678 241 2270 247
rect 2336 281 2928 287
rect 2336 247 2348 281
rect 2916 247 2928 281
rect 2336 241 2928 247
rect -2984 188 -2938 200
rect -2984 -188 -2978 188
rect -2944 -188 -2938 188
rect -2984 -200 -2938 -188
rect -2326 188 -2280 200
rect -2326 -188 -2320 188
rect -2286 -188 -2280 188
rect -2326 -200 -2280 -188
rect -1668 188 -1622 200
rect -1668 -188 -1662 188
rect -1628 -188 -1622 188
rect -1668 -200 -1622 -188
rect -1010 188 -964 200
rect -1010 -188 -1004 188
rect -970 -188 -964 188
rect -1010 -200 -964 -188
rect -352 188 -306 200
rect -352 -188 -346 188
rect -312 -188 -306 188
rect -352 -200 -306 -188
rect 306 188 352 200
rect 306 -188 312 188
rect 346 -188 352 188
rect 306 -200 352 -188
rect 964 188 1010 200
rect 964 -188 970 188
rect 1004 -188 1010 188
rect 964 -200 1010 -188
rect 1622 188 1668 200
rect 1622 -188 1628 188
rect 1662 -188 1668 188
rect 1622 -200 1668 -188
rect 2280 188 2326 200
rect 2280 -188 2286 188
rect 2320 -188 2326 188
rect 2280 -200 2326 -188
rect 2938 188 2984 200
rect 2938 -188 2944 188
rect 2978 -188 2984 188
rect 2938 -200 2984 -188
rect -2928 -247 -2336 -241
rect -2928 -281 -2916 -247
rect -2348 -281 -2336 -247
rect -2928 -287 -2336 -281
rect -2270 -247 -1678 -241
rect -2270 -281 -2258 -247
rect -1690 -281 -1678 -247
rect -2270 -287 -1678 -281
rect -1612 -247 -1020 -241
rect -1612 -281 -1600 -247
rect -1032 -281 -1020 -247
rect -1612 -287 -1020 -281
rect -954 -247 -362 -241
rect -954 -281 -942 -247
rect -374 -281 -362 -247
rect -954 -287 -362 -281
rect -296 -247 296 -241
rect -296 -281 -284 -247
rect 284 -281 296 -247
rect -296 -287 296 -281
rect 362 -247 954 -241
rect 362 -281 374 -247
rect 942 -281 954 -247
rect 362 -287 954 -281
rect 1020 -247 1612 -241
rect 1020 -281 1032 -247
rect 1600 -281 1612 -247
rect 1020 -287 1612 -281
rect 1678 -247 2270 -241
rect 1678 -281 1690 -247
rect 2258 -281 2270 -247
rect 1678 -287 2270 -281
rect 2336 -247 2928 -241
rect 2336 -281 2348 -247
rect 2916 -281 2928 -247
rect 2336 -287 2928 -281
<< properties >>
string FIXED_BBOX -3075 -366 3075 366
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 2.0 l 3.0 m 1 nf 9 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

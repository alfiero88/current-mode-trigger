magic
tech sky130A
magscale 1 2
timestamp 1716907293
<< error_p >>
rect -221 372 -163 378
rect -29 372 29 378
rect 163 372 221 378
rect -221 338 -209 372
rect -29 338 -17 372
rect 163 338 175 372
rect -221 332 -163 338
rect -29 332 29 338
rect 163 332 221 338
rect -317 -338 -259 -332
rect -125 -338 -67 -332
rect 67 -338 125 -332
rect 259 -338 317 -332
rect -317 -372 -305 -338
rect -125 -372 -113 -338
rect 67 -372 79 -338
rect 259 -372 271 -338
rect -317 -378 -259 -372
rect -125 -378 -67 -372
rect 67 -378 125 -372
rect 259 -378 317 -372
<< pwell >>
rect -503 -510 503 510
<< nmoslvt >>
rect -303 -300 -273 300
rect -207 -300 -177 300
rect -111 -300 -81 300
rect -15 -300 15 300
rect 81 -300 111 300
rect 177 -300 207 300
rect 273 -300 303 300
<< ndiff >>
rect -365 288 -303 300
rect -365 -288 -353 288
rect -319 -288 -303 288
rect -365 -300 -303 -288
rect -273 288 -207 300
rect -273 -288 -257 288
rect -223 -288 -207 288
rect -273 -300 -207 -288
rect -177 288 -111 300
rect -177 -288 -161 288
rect -127 -288 -111 288
rect -177 -300 -111 -288
rect -81 288 -15 300
rect -81 -288 -65 288
rect -31 -288 -15 288
rect -81 -300 -15 -288
rect 15 288 81 300
rect 15 -288 31 288
rect 65 -288 81 288
rect 15 -300 81 -288
rect 111 288 177 300
rect 111 -288 127 288
rect 161 -288 177 288
rect 111 -300 177 -288
rect 207 288 273 300
rect 207 -288 223 288
rect 257 -288 273 288
rect 207 -300 273 -288
rect 303 288 365 300
rect 303 -288 319 288
rect 353 -288 365 288
rect 303 -300 365 -288
<< ndiffc >>
rect -353 -288 -319 288
rect -257 -288 -223 288
rect -161 -288 -127 288
rect -65 -288 -31 288
rect 31 -288 65 288
rect 127 -288 161 288
rect 223 -288 257 288
rect 319 -288 353 288
<< psubdiff >>
rect -467 440 -371 474
rect 371 440 467 474
rect -467 378 -433 440
rect 433 378 467 440
rect -467 -440 -433 -378
rect 433 -440 467 -378
rect -467 -474 -371 -440
rect 371 -474 467 -440
<< psubdiffcont >>
rect -371 440 371 474
rect -467 -378 -433 378
rect 433 -378 467 378
rect -371 -474 371 -440
<< poly >>
rect -225 372 -159 388
rect -225 338 -209 372
rect -175 338 -159 372
rect -303 300 -273 326
rect -225 322 -159 338
rect -33 372 33 388
rect -33 338 -17 372
rect 17 338 33 372
rect -207 300 -177 322
rect -111 300 -81 326
rect -33 322 33 338
rect 159 372 225 388
rect 159 338 175 372
rect 209 338 225 372
rect -15 300 15 322
rect 81 300 111 326
rect 159 322 225 338
rect 177 300 207 322
rect 273 300 303 326
rect -303 -322 -273 -300
rect -321 -338 -255 -322
rect -207 -326 -177 -300
rect -111 -322 -81 -300
rect -321 -372 -305 -338
rect -271 -372 -255 -338
rect -321 -388 -255 -372
rect -129 -338 -63 -322
rect -15 -326 15 -300
rect 81 -322 111 -300
rect -129 -372 -113 -338
rect -79 -372 -63 -338
rect -129 -388 -63 -372
rect 63 -338 129 -322
rect 177 -326 207 -300
rect 273 -322 303 -300
rect 63 -372 79 -338
rect 113 -372 129 -338
rect 63 -388 129 -372
rect 255 -338 321 -322
rect 255 -372 271 -338
rect 305 -372 321 -338
rect 255 -388 321 -372
<< polycont >>
rect -209 338 -175 372
rect -17 338 17 372
rect 175 338 209 372
rect -305 -372 -271 -338
rect -113 -372 -79 -338
rect 79 -372 113 -338
rect 271 -372 305 -338
<< locali >>
rect -467 440 -371 474
rect 371 440 467 474
rect -467 378 -433 440
rect 433 378 467 440
rect -225 338 -209 372
rect -175 338 -159 372
rect -33 338 -17 372
rect 17 338 33 372
rect 159 338 175 372
rect 209 338 225 372
rect -353 288 -319 304
rect -353 -304 -319 -288
rect -257 288 -223 304
rect -257 -304 -223 -288
rect -161 288 -127 304
rect -161 -304 -127 -288
rect -65 288 -31 304
rect -65 -304 -31 -288
rect 31 288 65 304
rect 31 -304 65 -288
rect 127 288 161 304
rect 127 -304 161 -288
rect 223 288 257 304
rect 223 -304 257 -288
rect 319 288 353 304
rect 319 -304 353 -288
rect -321 -372 -305 -338
rect -271 -372 -255 -338
rect -129 -372 -113 -338
rect -79 -372 -63 -338
rect 63 -372 79 -338
rect 113 -372 129 -338
rect 255 -372 271 -338
rect 305 -372 321 -338
rect -467 -440 -433 -378
rect 433 -440 467 -378
rect -467 -474 -371 -440
rect 371 -474 467 -440
<< viali >>
rect -209 338 -175 372
rect -17 338 17 372
rect 175 338 209 372
rect -353 -288 -319 288
rect -257 -288 -223 288
rect -161 -288 -127 288
rect -65 -288 -31 288
rect 31 -288 65 288
rect 127 -288 161 288
rect 223 -288 257 288
rect 319 -288 353 288
rect -305 -372 -271 -338
rect -113 -372 -79 -338
rect 79 -372 113 -338
rect 271 -372 305 -338
<< metal1 >>
rect -221 372 -163 378
rect -221 338 -209 372
rect -175 338 -163 372
rect -221 332 -163 338
rect -29 372 29 378
rect -29 338 -17 372
rect 17 338 29 372
rect -29 332 29 338
rect 163 372 221 378
rect 163 338 175 372
rect 209 338 221 372
rect 163 332 221 338
rect -359 288 -313 300
rect -359 -288 -353 288
rect -319 -288 -313 288
rect -359 -300 -313 -288
rect -263 288 -217 300
rect -263 -288 -257 288
rect -223 -288 -217 288
rect -263 -300 -217 -288
rect -167 288 -121 300
rect -167 -288 -161 288
rect -127 -288 -121 288
rect -167 -300 -121 -288
rect -71 288 -25 300
rect -71 -288 -65 288
rect -31 -288 -25 288
rect -71 -300 -25 -288
rect 25 288 71 300
rect 25 -288 31 288
rect 65 -288 71 288
rect 25 -300 71 -288
rect 121 288 167 300
rect 121 -288 127 288
rect 161 -288 167 288
rect 121 -300 167 -288
rect 217 288 263 300
rect 217 -288 223 288
rect 257 -288 263 288
rect 217 -300 263 -288
rect 313 288 359 300
rect 313 -288 319 288
rect 353 -288 359 288
rect 313 -300 359 -288
rect -317 -338 -259 -332
rect -317 -372 -305 -338
rect -271 -372 -259 -338
rect -317 -378 -259 -372
rect -125 -338 -67 -332
rect -125 -372 -113 -338
rect -79 -372 -67 -338
rect -125 -378 -67 -372
rect 67 -338 125 -332
rect 67 -372 79 -338
rect 113 -372 125 -338
rect 67 -378 125 -372
rect 259 -338 317 -332
rect 259 -372 271 -338
rect 305 -372 317 -338
rect 259 -378 317 -372
<< properties >>
string FIXED_BBOX -450 -457 450 457
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 3.0 l 0.15 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
timestamp 1716907293
<< pwell >>
rect -277 -155 277 155
<< nmoslvt >>
rect -179 -50 -79 50
rect -50 -50 50 50
rect 79 -50 179 50
<< ndiff >>
rect -208 44 -179 50
rect -208 -44 -202 44
rect -185 -44 -179 44
rect -208 -50 -179 -44
rect -79 44 -50 50
rect -79 -44 -73 44
rect -56 -44 -50 44
rect -79 -50 -50 -44
rect 50 44 79 50
rect 50 -44 56 44
rect 73 -44 79 44
rect 50 -50 79 -44
rect 179 44 208 50
rect 179 -44 185 44
rect 202 -44 208 44
rect 179 -50 208 -44
<< ndiffc >>
rect -202 -44 -185 44
rect -73 -44 -56 44
rect 56 -44 73 44
rect 185 -44 202 44
<< psubdiff >>
rect -259 120 -211 137
rect 211 120 259 137
rect -259 89 -242 120
rect 242 89 259 120
rect -259 -120 -242 -89
rect 242 -120 259 -89
rect -259 -137 -211 -120
rect 211 -137 259 -120
<< psubdiffcont >>
rect -211 120 211 137
rect -259 -89 -242 89
rect 242 -89 259 89
rect -211 -137 211 -120
<< poly >>
rect -179 86 -79 94
rect -179 69 -171 86
rect -87 69 -79 86
rect -179 50 -79 69
rect -50 86 50 94
rect -50 69 -42 86
rect 42 69 50 86
rect -50 50 50 69
rect 79 86 179 94
rect 79 69 87 86
rect 171 69 179 86
rect 79 50 179 69
rect -179 -69 -79 -50
rect -179 -86 -171 -69
rect -87 -86 -79 -69
rect -179 -94 -79 -86
rect -50 -69 50 -50
rect -50 -86 -42 -69
rect 42 -86 50 -69
rect -50 -94 50 -86
rect 79 -69 179 -50
rect 79 -86 87 -69
rect 171 -86 179 -69
rect 79 -94 179 -86
<< polycont >>
rect -171 69 -87 86
rect -42 69 42 86
rect 87 69 171 86
rect -171 -86 -87 -69
rect -42 -86 42 -69
rect 87 -86 171 -69
<< locali >>
rect -259 120 -211 137
rect 211 120 259 137
rect -259 89 -242 120
rect 242 89 259 120
rect -179 69 -171 86
rect -87 69 -79 86
rect -50 69 -42 86
rect 42 69 50 86
rect 79 69 87 86
rect 171 69 179 86
rect -202 44 -185 52
rect -202 -52 -185 -44
rect -73 44 -56 52
rect -73 -52 -56 -44
rect 56 44 73 52
rect 56 -52 73 -44
rect 185 44 202 52
rect 185 -52 202 -44
rect -179 -86 -171 -69
rect -87 -86 -79 -69
rect -50 -86 -42 -69
rect 42 -86 50 -69
rect 79 -86 87 -69
rect 171 -86 179 -69
rect -259 -120 -242 -89
rect 242 -120 259 -89
rect -259 -137 -211 -120
rect 211 -137 259 -120
<< viali >>
rect -171 69 -87 86
rect -42 69 42 86
rect 87 69 171 86
rect -202 -44 -185 44
rect -73 -44 -56 44
rect 56 -44 73 44
rect 185 -44 202 44
rect -171 -86 -87 -69
rect -42 -86 42 -69
rect 87 -86 171 -69
<< metal1 >>
rect -177 86 -81 89
rect -177 69 -171 86
rect -87 69 -81 86
rect -177 66 -81 69
rect -48 86 48 89
rect -48 69 -42 86
rect 42 69 48 86
rect -48 66 48 69
rect 81 86 177 89
rect 81 69 87 86
rect 171 69 177 86
rect 81 66 177 69
rect -205 44 -182 50
rect -205 -44 -202 44
rect -185 -44 -182 44
rect -205 -50 -182 -44
rect -76 44 -53 50
rect -76 -44 -73 44
rect -56 -44 -53 44
rect -76 -50 -53 -44
rect 53 44 76 50
rect 53 -44 56 44
rect 73 -44 76 44
rect 53 -50 76 -44
rect 182 44 205 50
rect 182 -44 185 44
rect 202 -44 205 44
rect 182 -50 205 -44
rect -177 -69 -81 -66
rect -177 -86 -171 -69
rect -87 -86 -81 -69
rect -177 -89 -81 -86
rect -48 -69 48 -66
rect -48 -86 -42 -69
rect 42 -86 48 -69
rect -48 -89 48 -86
rect 81 -69 177 -66
rect 81 -86 87 -69
rect 171 -86 177 -69
rect 81 -89 177 -86
<< properties >>
string FIXED_BBOX -250 -128 250 128
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.0 l 1.0 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

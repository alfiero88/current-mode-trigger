magic
tech sky130A
magscale 1 2
timestamp 1717165854
<< metal1 >>
rect 25075 28838 29281 28956
rect 25075 28538 25192 28838
rect 25492 28538 29281 28838
rect 25075 28421 29281 28538
rect 19203 27322 21689 27425
rect 19203 27022 19306 27322
rect 19606 27022 21689 27322
rect 19203 26919 21689 27022
rect 21183 25347 21689 26919
rect 25300 26650 27487 26709
rect 25300 26470 27248 26650
rect 27428 26470 27487 26650
rect 25300 26412 27487 26470
rect 25300 25568 25597 26412
rect 28746 25215 29281 28421
rect 22218 13850 23354 13906
rect 22218 13670 22274 13850
rect 22454 13670 23354 13850
rect 22218 13614 23354 13670
rect 26607 7072 26849 7859
rect 26607 6892 26638 7072
rect 26818 6892 26849 7072
rect 26607 6861 26849 6892
rect 24579 5328 24861 6397
rect 24579 5148 24630 5328
rect 24810 5148 24861 5328
rect 24579 5097 24861 5148
<< via1 >>
rect 25192 28538 25492 28838
rect 19306 27022 19606 27322
rect 27248 26470 27428 26650
rect 22274 13670 22454 13850
rect 26638 6892 26818 7072
rect 24630 5148 24810 5328
<< metal2 >>
rect 17445 28838 17735 28842
rect 17440 28833 25192 28838
rect 17440 28543 17445 28833
rect 17735 28543 25192 28833
rect 17440 28538 25192 28543
rect 25492 28538 25498 28838
rect 17445 28534 17735 28538
rect 17387 27322 17677 27326
rect 17382 27317 19306 27322
rect 17382 27027 17387 27317
rect 17677 27027 19306 27317
rect 17382 27022 19306 27027
rect 19606 27022 19612 27322
rect 17387 27018 17677 27022
rect 27242 26470 27248 26650
rect 27428 26470 31462 26650
rect 31282 23211 31462 26470
rect 31278 23041 31287 23211
rect 31457 23041 31466 23211
rect 31282 23036 31462 23041
rect 18034 13670 22274 13850
rect 22454 13670 22460 13850
rect 18034 12857 18214 13670
rect 18030 12687 18039 12857
rect 18209 12687 18218 12857
rect 18034 12682 18214 12687
rect 26638 7072 26818 7078
rect 24630 5328 24810 5334
rect 24630 4245 24810 5148
rect 26638 4391 26818 6892
rect 24626 4075 24635 4245
rect 24805 4075 24814 4245
rect 26634 4221 26643 4391
rect 26813 4221 26822 4391
rect 26638 4216 26818 4221
rect 24630 4070 24810 4075
<< via2 >>
rect 17445 28543 17735 28833
rect 17387 27027 17677 27317
rect 31287 23041 31457 23211
rect 18039 12687 18209 12857
rect 24635 4075 24805 4245
rect 26643 4221 26813 4391
<< metal3 >>
rect 5785 28838 6083 28843
rect 5784 28837 17740 28838
rect 5784 28539 5785 28837
rect 6083 28833 17740 28837
rect 6083 28543 17445 28833
rect 17735 28543 17740 28833
rect 6083 28539 17740 28543
rect 5784 28538 17740 28539
rect 5785 28533 6083 28538
rect 15693 27322 15991 27327
rect 15692 27321 17682 27322
rect 15692 27023 15693 27321
rect 15991 27317 17682 27321
rect 15991 27027 17387 27317
rect 17677 27027 17682 27317
rect 15991 27023 17682 27027
rect 15692 27022 17682 27023
rect 15693 27017 15991 27022
rect 31282 23211 31462 23216
rect 31282 23041 31287 23211
rect 31457 23041 31462 23211
rect 31282 14023 31462 23041
rect 31282 13845 31283 14023
rect 31461 13845 31462 14023
rect 31282 13844 31462 13845
rect 31283 13839 31461 13844
rect 18034 12857 18214 12862
rect 18034 12687 18039 12857
rect 18209 12687 18214 12857
rect 18034 7449 18214 12687
rect 18029 7271 18035 7449
rect 18213 7271 18219 7449
rect 18034 7270 18214 7271
rect 26638 4391 26818 4396
rect 24630 4245 24810 4250
rect 24630 4075 24635 4245
rect 24805 4075 24810 4245
rect 24630 2795 24810 4075
rect 26638 4221 26643 4391
rect 26813 4221 26818 4391
rect 26638 3087 26818 4221
rect 26633 2909 26639 3087
rect 26817 2909 26823 3087
rect 26638 2908 26818 2909
rect 24625 2617 24631 2795
rect 24809 2617 24815 2795
rect 24630 2616 24810 2617
<< via3 >>
rect 5785 28539 6083 28837
rect 15693 27023 15991 27321
rect 31283 13845 31461 14023
rect 18035 7271 18213 7449
rect 26639 2909 26817 3087
rect 24631 2617 24809 2795
<< metal4 >>
rect 798 44822 858 45152
rect 1534 44822 1594 45152
rect 2270 44822 2330 45152
rect 3006 44822 3066 45152
rect 3742 44822 3802 45152
rect 4478 44822 4538 45152
rect 5214 44822 5274 45152
rect 5950 44822 6010 45152
rect 6686 44822 6746 45152
rect 7422 44822 7482 45152
rect 8158 44822 8218 45152
rect 8894 44822 8954 45152
rect 9630 44822 9690 45152
rect 10366 44822 10426 45152
rect 11102 44822 11162 45152
rect 11838 44822 11898 45152
rect 12574 44822 12634 45152
rect 13310 44822 13370 45152
rect 14046 44822 14106 45152
rect 14782 44822 14842 45152
rect 15518 44822 15578 45152
rect 16254 44822 16314 45152
rect 16990 44822 17050 45152
rect 17726 44822 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 620 44528 17852 44822
rect 200 28838 500 44152
rect 200 28837 6084 28838
rect 200 28539 5785 28837
rect 6083 28539 6084 28837
rect 200 28538 6084 28539
rect 200 1000 500 28538
rect 9800 27322 10100 44528
rect 9800 27321 15992 27322
rect 9800 27023 15693 27321
rect 15991 27023 15992 27321
rect 9800 27022 15992 27023
rect 9800 1000 10100 27022
rect 31282 14023 31462 14024
rect 31282 13845 31283 14023
rect 31461 13845 31462 14023
rect 18034 7449 18214 7450
rect 18034 7271 18035 7449
rect 18213 7271 18214 7449
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 7271
rect 26638 3087 26818 3088
rect 26638 2909 26639 3087
rect 26817 2909 26818 3087
rect 24630 2795 24810 2796
rect 24630 2617 24631 2795
rect 24809 2617 24810 2795
rect 24630 1372 24810 2617
rect 26638 2040 26818 2909
rect 26638 1860 27046 2040
rect 22450 1192 24810 1372
rect 22450 0 22630 1192
rect 26866 0 27046 1860
rect 31282 0 31462 13845
use CurrentTrigger  CurrentTrigger_0
timestamp 1717084777
transform 0 1 19364 -1 0 25020
box -854 1682 19074 10100
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 4800 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 4800 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>

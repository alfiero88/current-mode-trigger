magic
tech sky130A
magscale 1 2
timestamp 1716907293
<< nwell >>
rect -2141 -419 2141 419
<< pmoslvt >>
rect -1945 -200 -1345 200
rect -1287 -200 -687 200
rect -629 -200 -29 200
rect 29 -200 629 200
rect 687 -200 1287 200
rect 1345 -200 1945 200
<< pdiff >>
rect -2003 188 -1945 200
rect -2003 -188 -1991 188
rect -1957 -188 -1945 188
rect -2003 -200 -1945 -188
rect -1345 188 -1287 200
rect -1345 -188 -1333 188
rect -1299 -188 -1287 188
rect -1345 -200 -1287 -188
rect -687 188 -629 200
rect -687 -188 -675 188
rect -641 -188 -629 188
rect -687 -200 -629 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 629 188 687 200
rect 629 -188 641 188
rect 675 -188 687 188
rect 629 -200 687 -188
rect 1287 188 1345 200
rect 1287 -188 1299 188
rect 1333 -188 1345 188
rect 1287 -200 1345 -188
rect 1945 188 2003 200
rect 1945 -188 1957 188
rect 1991 -188 2003 188
rect 1945 -200 2003 -188
<< pdiffc >>
rect -1991 -188 -1957 188
rect -1333 -188 -1299 188
rect -675 -188 -641 188
rect -17 -188 17 188
rect 641 -188 675 188
rect 1299 -188 1333 188
rect 1957 -188 1991 188
<< nsubdiff >>
rect -2105 349 -2009 383
rect 2009 349 2105 383
rect -2105 287 -2071 349
rect 2071 287 2105 349
rect -2105 -349 -2071 -287
rect 2071 -349 2105 -287
rect -2105 -383 -2009 -349
rect 2009 -383 2105 -349
<< nsubdiffcont >>
rect -2009 349 2009 383
rect -2105 -287 -2071 287
rect 2071 -287 2105 287
rect -2009 -383 2009 -349
<< poly >>
rect -1945 281 -1345 297
rect -1945 247 -1929 281
rect -1361 247 -1345 281
rect -1945 200 -1345 247
rect -1287 281 -687 297
rect -1287 247 -1271 281
rect -703 247 -687 281
rect -1287 200 -687 247
rect -629 281 -29 297
rect -629 247 -613 281
rect -45 247 -29 281
rect -629 200 -29 247
rect 29 281 629 297
rect 29 247 45 281
rect 613 247 629 281
rect 29 200 629 247
rect 687 281 1287 297
rect 687 247 703 281
rect 1271 247 1287 281
rect 687 200 1287 247
rect 1345 281 1945 297
rect 1345 247 1361 281
rect 1929 247 1945 281
rect 1345 200 1945 247
rect -1945 -247 -1345 -200
rect -1945 -281 -1929 -247
rect -1361 -281 -1345 -247
rect -1945 -297 -1345 -281
rect -1287 -247 -687 -200
rect -1287 -281 -1271 -247
rect -703 -281 -687 -247
rect -1287 -297 -687 -281
rect -629 -247 -29 -200
rect -629 -281 -613 -247
rect -45 -281 -29 -247
rect -629 -297 -29 -281
rect 29 -247 629 -200
rect 29 -281 45 -247
rect 613 -281 629 -247
rect 29 -297 629 -281
rect 687 -247 1287 -200
rect 687 -281 703 -247
rect 1271 -281 1287 -247
rect 687 -297 1287 -281
rect 1345 -247 1945 -200
rect 1345 -281 1361 -247
rect 1929 -281 1945 -247
rect 1345 -297 1945 -281
<< polycont >>
rect -1929 247 -1361 281
rect -1271 247 -703 281
rect -613 247 -45 281
rect 45 247 613 281
rect 703 247 1271 281
rect 1361 247 1929 281
rect -1929 -281 -1361 -247
rect -1271 -281 -703 -247
rect -613 -281 -45 -247
rect 45 -281 613 -247
rect 703 -281 1271 -247
rect 1361 -281 1929 -247
<< locali >>
rect -2105 349 -2009 383
rect 2009 349 2105 383
rect -2105 287 -2071 349
rect 2071 287 2105 349
rect -1945 247 -1929 281
rect -1361 247 -1345 281
rect -1287 247 -1271 281
rect -703 247 -687 281
rect -629 247 -613 281
rect -45 247 -29 281
rect 29 247 45 281
rect 613 247 629 281
rect 687 247 703 281
rect 1271 247 1287 281
rect 1345 247 1361 281
rect 1929 247 1945 281
rect -1991 188 -1957 204
rect -1991 -204 -1957 -188
rect -1333 188 -1299 204
rect -1333 -204 -1299 -188
rect -675 188 -641 204
rect -675 -204 -641 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 641 188 675 204
rect 641 -204 675 -188
rect 1299 188 1333 204
rect 1299 -204 1333 -188
rect 1957 188 1991 204
rect 1957 -204 1991 -188
rect -1945 -281 -1929 -247
rect -1361 -281 -1345 -247
rect -1287 -281 -1271 -247
rect -703 -281 -687 -247
rect -629 -281 -613 -247
rect -45 -281 -29 -247
rect 29 -281 45 -247
rect 613 -281 629 -247
rect 687 -281 703 -247
rect 1271 -281 1287 -247
rect 1345 -281 1361 -247
rect 1929 -281 1945 -247
rect -2105 -349 -2071 -287
rect 2071 -349 2105 -287
rect -2105 -383 -2009 -349
rect 2009 -383 2105 -349
<< viali >>
rect -1929 247 -1361 281
rect -1271 247 -703 281
rect -613 247 -45 281
rect 45 247 613 281
rect 703 247 1271 281
rect 1361 247 1929 281
rect -1991 -188 -1957 188
rect -1333 -188 -1299 188
rect -675 -188 -641 188
rect -17 -188 17 188
rect 641 -188 675 188
rect 1299 -188 1333 188
rect 1957 -188 1991 188
rect -1929 -281 -1361 -247
rect -1271 -281 -703 -247
rect -613 -281 -45 -247
rect 45 -281 613 -247
rect 703 -281 1271 -247
rect 1361 -281 1929 -247
<< metal1 >>
rect -1941 281 -1349 287
rect -1941 247 -1929 281
rect -1361 247 -1349 281
rect -1941 241 -1349 247
rect -1283 281 -691 287
rect -1283 247 -1271 281
rect -703 247 -691 281
rect -1283 241 -691 247
rect -625 281 -33 287
rect -625 247 -613 281
rect -45 247 -33 281
rect -625 241 -33 247
rect 33 281 625 287
rect 33 247 45 281
rect 613 247 625 281
rect 33 241 625 247
rect 691 281 1283 287
rect 691 247 703 281
rect 1271 247 1283 281
rect 691 241 1283 247
rect 1349 281 1941 287
rect 1349 247 1361 281
rect 1929 247 1941 281
rect 1349 241 1941 247
rect -1997 188 -1951 200
rect -1997 -188 -1991 188
rect -1957 -188 -1951 188
rect -1997 -200 -1951 -188
rect -1339 188 -1293 200
rect -1339 -188 -1333 188
rect -1299 -188 -1293 188
rect -1339 -200 -1293 -188
rect -681 188 -635 200
rect -681 -188 -675 188
rect -641 -188 -635 188
rect -681 -200 -635 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 635 188 681 200
rect 635 -188 641 188
rect 675 -188 681 188
rect 635 -200 681 -188
rect 1293 188 1339 200
rect 1293 -188 1299 188
rect 1333 -188 1339 188
rect 1293 -200 1339 -188
rect 1951 188 1997 200
rect 1951 -188 1957 188
rect 1991 -188 1997 188
rect 1951 -200 1997 -188
rect -1941 -247 -1349 -241
rect -1941 -281 -1929 -247
rect -1361 -281 -1349 -247
rect -1941 -287 -1349 -281
rect -1283 -247 -691 -241
rect -1283 -281 -1271 -247
rect -703 -281 -691 -247
rect -1283 -287 -691 -281
rect -625 -247 -33 -241
rect -625 -281 -613 -247
rect -45 -281 -33 -247
rect -625 -287 -33 -281
rect 33 -247 625 -241
rect 33 -281 45 -247
rect 613 -281 625 -247
rect 33 -287 625 -281
rect 691 -247 1283 -241
rect 691 -281 703 -247
rect 1271 -281 1283 -247
rect 691 -287 1283 -281
rect 1349 -247 1941 -241
rect 1349 -281 1361 -247
rect 1929 -281 1941 -247
rect 1349 -287 1941 -281
<< properties >>
string FIXED_BBOX -2088 -366 2088 366
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 2.0 l 3.0 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

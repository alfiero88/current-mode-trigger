magic
tech sky130A
magscale 1 2
timestamp 1716907293
<< error_p >>
rect -415 295 -353 301
rect -287 295 -225 301
rect -159 295 -97 301
rect -31 295 31 301
rect 97 295 159 301
rect 225 295 287 301
rect 353 295 415 301
rect -415 261 -403 295
rect -287 261 -275 295
rect -159 261 -147 295
rect -31 261 -19 295
rect 97 261 109 295
rect 225 261 237 295
rect 353 261 365 295
rect -415 255 -353 261
rect -287 255 -225 261
rect -159 255 -97 261
rect -31 255 31 261
rect 97 255 159 261
rect 225 255 287 261
rect 353 255 415 261
rect -415 -261 -353 -255
rect -287 -261 -225 -255
rect -159 -261 -97 -255
rect -31 -261 31 -255
rect 97 -261 159 -255
rect 225 -261 287 -255
rect 353 -261 415 -255
rect -415 -295 -403 -261
rect -287 -295 -275 -261
rect -159 -295 -147 -261
rect -31 -295 -19 -261
rect 97 -295 109 -261
rect 225 -295 237 -261
rect 353 -295 365 -261
rect -415 -301 -353 -295
rect -287 -301 -225 -295
rect -159 -301 -97 -295
rect -31 -301 31 -295
rect 97 -301 159 -295
rect 225 -301 287 -295
rect 353 -301 415 -295
<< nwell >>
rect -615 -433 615 433
<< pmoslvt >>
rect -419 -214 -349 214
rect -291 -214 -221 214
rect -163 -214 -93 214
rect -35 -214 35 214
rect 93 -214 163 214
rect 221 -214 291 214
rect 349 -214 419 214
<< pdiff >>
rect -477 202 -419 214
rect -477 -202 -465 202
rect -431 -202 -419 202
rect -477 -214 -419 -202
rect -349 202 -291 214
rect -349 -202 -337 202
rect -303 -202 -291 202
rect -349 -214 -291 -202
rect -221 202 -163 214
rect -221 -202 -209 202
rect -175 -202 -163 202
rect -221 -214 -163 -202
rect -93 202 -35 214
rect -93 -202 -81 202
rect -47 -202 -35 202
rect -93 -214 -35 -202
rect 35 202 93 214
rect 35 -202 47 202
rect 81 -202 93 202
rect 35 -214 93 -202
rect 163 202 221 214
rect 163 -202 175 202
rect 209 -202 221 202
rect 163 -214 221 -202
rect 291 202 349 214
rect 291 -202 303 202
rect 337 -202 349 202
rect 291 -214 349 -202
rect 419 202 477 214
rect 419 -202 431 202
rect 465 -202 477 202
rect 419 -214 477 -202
<< pdiffc >>
rect -465 -202 -431 202
rect -337 -202 -303 202
rect -209 -202 -175 202
rect -81 -202 -47 202
rect 47 -202 81 202
rect 175 -202 209 202
rect 303 -202 337 202
rect 431 -202 465 202
<< nsubdiff >>
rect -579 363 -483 397
rect 483 363 579 397
rect -579 301 -545 363
rect 545 301 579 363
rect -579 -363 -545 -301
rect 545 -363 579 -301
rect -579 -397 -483 -363
rect 483 -397 579 -363
<< nsubdiffcont >>
rect -483 363 483 397
rect -579 -301 -545 301
rect 545 -301 579 301
rect -483 -397 483 -363
<< poly >>
rect -419 295 -349 311
rect -419 261 -403 295
rect -365 261 -349 295
rect -419 214 -349 261
rect -291 295 -221 311
rect -291 261 -275 295
rect -237 261 -221 295
rect -291 214 -221 261
rect -163 295 -93 311
rect -163 261 -147 295
rect -109 261 -93 295
rect -163 214 -93 261
rect -35 295 35 311
rect -35 261 -19 295
rect 19 261 35 295
rect -35 214 35 261
rect 93 295 163 311
rect 93 261 109 295
rect 147 261 163 295
rect 93 214 163 261
rect 221 295 291 311
rect 221 261 237 295
rect 275 261 291 295
rect 221 214 291 261
rect 349 295 419 311
rect 349 261 365 295
rect 403 261 419 295
rect 349 214 419 261
rect -419 -261 -349 -214
rect -419 -295 -403 -261
rect -365 -295 -349 -261
rect -419 -311 -349 -295
rect -291 -261 -221 -214
rect -291 -295 -275 -261
rect -237 -295 -221 -261
rect -291 -311 -221 -295
rect -163 -261 -93 -214
rect -163 -295 -147 -261
rect -109 -295 -93 -261
rect -163 -311 -93 -295
rect -35 -261 35 -214
rect -35 -295 -19 -261
rect 19 -295 35 -261
rect -35 -311 35 -295
rect 93 -261 163 -214
rect 93 -295 109 -261
rect 147 -295 163 -261
rect 93 -311 163 -295
rect 221 -261 291 -214
rect 221 -295 237 -261
rect 275 -295 291 -261
rect 221 -311 291 -295
rect 349 -261 419 -214
rect 349 -295 365 -261
rect 403 -295 419 -261
rect 349 -311 419 -295
<< polycont >>
rect -403 261 -365 295
rect -275 261 -237 295
rect -147 261 -109 295
rect -19 261 19 295
rect 109 261 147 295
rect 237 261 275 295
rect 365 261 403 295
rect -403 -295 -365 -261
rect -275 -295 -237 -261
rect -147 -295 -109 -261
rect -19 -295 19 -261
rect 109 -295 147 -261
rect 237 -295 275 -261
rect 365 -295 403 -261
<< locali >>
rect -579 363 -483 397
rect 483 363 579 397
rect -579 301 -545 363
rect 545 301 579 363
rect -419 261 -403 295
rect -365 261 -349 295
rect -291 261 -275 295
rect -237 261 -221 295
rect -163 261 -147 295
rect -109 261 -93 295
rect -35 261 -19 295
rect 19 261 35 295
rect 93 261 109 295
rect 147 261 163 295
rect 221 261 237 295
rect 275 261 291 295
rect 349 261 365 295
rect 403 261 419 295
rect -465 202 -431 218
rect -465 -218 -431 -202
rect -337 202 -303 218
rect -337 -218 -303 -202
rect -209 202 -175 218
rect -209 -218 -175 -202
rect -81 202 -47 218
rect -81 -218 -47 -202
rect 47 202 81 218
rect 47 -218 81 -202
rect 175 202 209 218
rect 175 -218 209 -202
rect 303 202 337 218
rect 303 -218 337 -202
rect 431 202 465 218
rect 431 -218 465 -202
rect -419 -295 -403 -261
rect -365 -295 -349 -261
rect -291 -295 -275 -261
rect -237 -295 -221 -261
rect -163 -295 -147 -261
rect -109 -295 -93 -261
rect -35 -295 -19 -261
rect 19 -295 35 -261
rect 93 -295 109 -261
rect 147 -295 163 -261
rect 221 -295 237 -261
rect 275 -295 291 -261
rect 349 -295 365 -261
rect 403 -295 419 -261
rect -579 -363 -545 -301
rect 545 -363 579 -301
rect -579 -397 -483 -363
rect 483 -397 579 -363
<< viali >>
rect -403 261 -365 295
rect -275 261 -237 295
rect -147 261 -109 295
rect -19 261 19 295
rect 109 261 147 295
rect 237 261 275 295
rect 365 261 403 295
rect -465 -202 -431 202
rect -337 -202 -303 202
rect -209 -202 -175 202
rect -81 -202 -47 202
rect 47 -202 81 202
rect 175 -202 209 202
rect 303 -202 337 202
rect 431 -202 465 202
rect -403 -295 -365 -261
rect -275 -295 -237 -261
rect -147 -295 -109 -261
rect -19 -295 19 -261
rect 109 -295 147 -261
rect 237 -295 275 -261
rect 365 -295 403 -261
<< metal1 >>
rect -415 295 -353 301
rect -415 261 -403 295
rect -365 261 -353 295
rect -415 255 -353 261
rect -287 295 -225 301
rect -287 261 -275 295
rect -237 261 -225 295
rect -287 255 -225 261
rect -159 295 -97 301
rect -159 261 -147 295
rect -109 261 -97 295
rect -159 255 -97 261
rect -31 295 31 301
rect -31 261 -19 295
rect 19 261 31 295
rect -31 255 31 261
rect 97 295 159 301
rect 97 261 109 295
rect 147 261 159 295
rect 97 255 159 261
rect 225 295 287 301
rect 225 261 237 295
rect 275 261 287 295
rect 225 255 287 261
rect 353 295 415 301
rect 353 261 365 295
rect 403 261 415 295
rect 353 255 415 261
rect -471 202 -425 214
rect -471 -202 -465 202
rect -431 -202 -425 202
rect -471 -214 -425 -202
rect -343 202 -297 214
rect -343 -202 -337 202
rect -303 -202 -297 202
rect -343 -214 -297 -202
rect -215 202 -169 214
rect -215 -202 -209 202
rect -175 -202 -169 202
rect -215 -214 -169 -202
rect -87 202 -41 214
rect -87 -202 -81 202
rect -47 -202 -41 202
rect -87 -214 -41 -202
rect 41 202 87 214
rect 41 -202 47 202
rect 81 -202 87 202
rect 41 -214 87 -202
rect 169 202 215 214
rect 169 -202 175 202
rect 209 -202 215 202
rect 169 -214 215 -202
rect 297 202 343 214
rect 297 -202 303 202
rect 337 -202 343 202
rect 297 -214 343 -202
rect 425 202 471 214
rect 425 -202 431 202
rect 465 -202 471 202
rect 425 -214 471 -202
rect -415 -261 -353 -255
rect -415 -295 -403 -261
rect -365 -295 -353 -261
rect -415 -301 -353 -295
rect -287 -261 -225 -255
rect -287 -295 -275 -261
rect -237 -295 -225 -261
rect -287 -301 -225 -295
rect -159 -261 -97 -255
rect -159 -295 -147 -261
rect -109 -295 -97 -261
rect -159 -301 -97 -295
rect -31 -261 31 -255
rect -31 -295 -19 -261
rect 19 -295 31 -261
rect -31 -301 31 -295
rect 97 -261 159 -255
rect 97 -295 109 -261
rect 147 -295 159 -261
rect 97 -301 159 -295
rect 225 -261 287 -255
rect 225 -295 237 -261
rect 275 -295 287 -261
rect 225 -301 287 -295
rect 353 -261 415 -255
rect 353 -295 365 -261
rect 403 -295 415 -261
rect 353 -301 415 -295
<< properties >>
string FIXED_BBOX -562 -380 562 380
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 2.142857142857143 l 0.35 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

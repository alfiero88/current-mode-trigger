VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_alfiero88_CurrentTrigger
  CLASS BLOCK ;
  FOREIGN tt_um_alfiero88_CurrentTrigger ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.350000 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.000000 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.530000 ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 10.312400 ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 111.090 114.940 116.190 119.900 ;
        RECT 120.750 114.870 125.850 119.900 ;
      LAYER nwell ;
        RECT 129.880 113.750 135.070 119.900 ;
        RECT 138.270 114.830 143.460 119.790 ;
      LAYER pwell ;
        RECT 111.670 93.190 117.770 104.730 ;
        RECT 111.730 77.590 117.830 89.130 ;
      LAYER nwell ;
        RECT 122.500 81.590 126.190 101.080 ;
        RECT 130.330 81.590 134.020 101.080 ;
      LAYER pwell ;
        RECT 114.720 68.440 117.820 73.980 ;
      LAYER nwell ;
        RECT 127.860 68.340 132.190 74.490 ;
        RECT 138.170 66.430 142.360 97.710 ;
      LAYER pwell ;
        RECT 114.750 54.470 117.850 60.010 ;
        RECT 128.990 52.920 132.090 61.460 ;
      LAYER nwell ;
        RECT 137.820 57.040 141.680 60.630 ;
      LAYER pwell ;
        RECT 120.520 44.480 123.620 46.590 ;
      LAYER nwell ;
        RECT 125.850 44.330 130.040 46.640 ;
      LAYER pwell ;
        RECT 120.520 39.280 124.120 41.910 ;
      LAYER nwell ;
        RECT 125.850 38.910 130.040 42.500 ;
      LAYER pwell ;
        RECT 119.080 31.970 124.180 35.080 ;
      LAYER nwell ;
        RECT 125.850 30.770 131.040 36.280 ;
        RECT 137.620 30.660 141.810 52.070 ;
      LAYER li1 ;
        RECT 121.380 119.720 125.230 119.770 ;
        RECT 130.520 119.720 134.420 119.750 ;
        RECT 111.270 119.550 116.010 119.720 ;
        RECT 111.270 119.270 111.440 119.550 ;
        RECT 111.230 115.580 111.440 119.270 ;
        RECT 112.120 118.980 115.160 119.150 ;
        RECT 111.780 115.920 111.950 118.920 ;
        RECT 115.330 115.920 115.500 118.920 ;
        RECT 112.120 115.690 115.160 115.860 ;
        RECT 111.270 115.290 111.440 115.580 ;
        RECT 115.840 115.290 116.010 119.550 ;
        RECT 111.270 115.120 116.010 115.290 ;
        RECT 120.930 119.550 125.670 119.720 ;
        RECT 120.930 115.220 121.100 119.550 ;
        RECT 121.440 118.660 121.610 118.990 ;
        RECT 121.780 118.980 124.820 119.150 ;
        RECT 121.780 118.500 124.820 118.670 ;
        RECT 121.440 117.700 121.610 118.030 ;
        RECT 121.780 118.020 124.820 118.190 ;
        RECT 124.990 118.180 125.160 118.510 ;
        RECT 121.780 117.540 124.820 117.710 ;
        RECT 121.440 116.740 121.610 117.070 ;
        RECT 121.780 117.060 124.820 117.230 ;
        RECT 124.990 117.220 125.160 117.550 ;
        RECT 121.780 116.580 124.820 116.750 ;
        RECT 121.440 115.780 121.610 116.110 ;
        RECT 121.780 116.100 124.820 116.270 ;
        RECT 124.990 116.260 125.160 116.590 ;
        RECT 121.780 115.620 124.820 115.790 ;
        RECT 125.500 115.220 125.670 119.550 ;
        RECT 120.930 115.050 125.670 115.220 ;
        RECT 130.060 119.550 134.890 119.720 ;
        RECT 130.060 114.100 130.230 119.550 ;
        RECT 130.955 118.980 133.995 119.150 ;
        RECT 130.570 118.570 130.740 118.920 ;
        RECT 134.210 118.570 134.380 118.920 ;
        RECT 130.955 118.340 133.995 118.510 ;
        RECT 130.570 117.930 130.740 118.280 ;
        RECT 134.210 117.930 134.380 118.280 ;
        RECT 130.955 117.700 133.995 117.870 ;
        RECT 130.570 117.290 130.740 117.640 ;
        RECT 134.210 117.290 134.380 117.640 ;
        RECT 130.955 117.060 133.995 117.230 ;
        RECT 130.570 116.650 130.740 117.000 ;
        RECT 134.210 116.650 134.380 117.000 ;
        RECT 130.955 116.420 133.995 116.590 ;
        RECT 130.570 116.010 130.740 116.360 ;
        RECT 134.210 116.010 134.380 116.360 ;
        RECT 130.955 115.780 133.995 115.950 ;
        RECT 130.570 115.370 130.740 115.720 ;
        RECT 134.210 115.370 134.380 115.720 ;
        RECT 130.955 115.140 133.995 115.310 ;
        RECT 130.570 114.730 130.740 115.080 ;
        RECT 134.210 114.730 134.380 115.080 ;
        RECT 130.955 114.500 133.995 114.670 ;
        RECT 134.720 114.100 134.890 119.550 ;
        RECT 138.450 119.440 143.280 119.610 ;
        RECT 138.450 115.180 138.620 119.440 ;
        RECT 143.110 119.150 143.280 119.440 ;
        RECT 139.345 118.870 142.385 119.040 ;
        RECT 138.960 115.810 139.130 118.810 ;
        RECT 142.600 115.810 142.770 118.810 ;
        RECT 139.345 115.580 142.385 115.750 ;
        RECT 143.110 115.470 143.310 119.150 ;
        RECT 143.110 115.180 143.280 115.470 ;
        RECT 138.450 115.010 143.280 115.180 ;
        RECT 130.060 113.930 134.890 114.100 ;
        RECT 111.850 104.380 117.590 104.550 ;
        RECT 111.850 104.100 112.020 104.380 ;
        RECT 111.780 93.820 112.020 104.100 ;
        RECT 112.700 103.810 116.740 103.980 ;
        RECT 112.360 100.750 112.530 103.750 ;
        RECT 116.910 100.750 117.080 103.750 ;
        RECT 112.700 100.520 116.740 100.690 ;
        RECT 112.360 97.460 112.530 100.460 ;
        RECT 116.910 97.460 117.080 100.460 ;
        RECT 112.700 97.230 116.740 97.400 ;
        RECT 112.360 94.170 112.530 97.170 ;
        RECT 116.910 94.170 117.080 97.170 ;
        RECT 112.700 93.940 116.740 94.110 ;
        RECT 111.850 93.540 112.020 93.820 ;
        RECT 117.420 93.540 117.590 104.380 ;
        RECT 111.850 93.370 117.590 93.540 ;
        RECT 122.680 100.730 126.010 100.900 ;
        RECT 111.910 88.780 117.650 88.950 ;
        RECT 111.910 88.490 112.080 88.780 ;
        RECT 111.840 78.230 112.080 88.490 ;
        RECT 112.760 88.210 116.800 88.380 ;
        RECT 112.420 85.150 112.590 88.150 ;
        RECT 116.970 85.150 117.140 88.150 ;
        RECT 112.760 84.920 116.800 85.090 ;
        RECT 112.420 81.860 112.590 84.860 ;
        RECT 116.970 81.860 117.140 84.860 ;
        RECT 112.760 81.630 116.800 81.800 ;
        RECT 112.420 78.570 112.590 81.570 ;
        RECT 116.970 78.570 117.140 81.570 ;
        RECT 112.760 78.340 116.800 78.510 ;
        RECT 111.910 77.940 112.080 78.230 ;
        RECT 117.480 77.940 117.650 88.780 ;
        RECT 122.680 81.940 122.850 100.730 ;
        RECT 125.840 100.470 126.010 100.730 ;
        RECT 130.510 100.730 133.840 100.900 ;
        RECT 123.575 100.160 125.115 100.330 ;
        RECT 123.190 99.400 123.360 100.100 ;
        RECT 125.330 99.400 125.500 100.100 ;
        RECT 123.575 99.170 125.115 99.340 ;
        RECT 123.190 98.410 123.360 99.110 ;
        RECT 125.330 98.410 125.500 99.110 ;
        RECT 123.575 98.180 125.115 98.350 ;
        RECT 123.190 97.420 123.360 98.120 ;
        RECT 125.330 97.420 125.500 98.120 ;
        RECT 123.575 97.190 125.115 97.360 ;
        RECT 123.190 96.430 123.360 97.130 ;
        RECT 125.330 96.430 125.500 97.130 ;
        RECT 123.575 96.200 125.115 96.370 ;
        RECT 123.190 95.440 123.360 96.140 ;
        RECT 125.330 95.440 125.500 96.140 ;
        RECT 123.575 95.210 125.115 95.380 ;
        RECT 123.190 94.450 123.360 95.150 ;
        RECT 125.330 94.450 125.500 95.150 ;
        RECT 123.575 94.220 125.115 94.390 ;
        RECT 123.190 93.460 123.360 94.160 ;
        RECT 125.330 93.460 125.500 94.160 ;
        RECT 123.575 93.230 125.115 93.400 ;
        RECT 123.190 92.470 123.360 93.170 ;
        RECT 125.330 92.470 125.500 93.170 ;
        RECT 123.575 92.240 125.115 92.410 ;
        RECT 123.190 91.480 123.360 92.180 ;
        RECT 125.330 91.480 125.500 92.180 ;
        RECT 123.575 91.250 125.115 91.420 ;
        RECT 123.190 90.490 123.360 91.190 ;
        RECT 125.330 90.490 125.500 91.190 ;
        RECT 123.575 90.260 125.115 90.430 ;
        RECT 123.190 89.500 123.360 90.200 ;
        RECT 125.330 89.500 125.500 90.200 ;
        RECT 123.575 89.270 125.115 89.440 ;
        RECT 123.190 88.510 123.360 89.210 ;
        RECT 125.330 88.510 125.500 89.210 ;
        RECT 123.575 88.280 125.115 88.450 ;
        RECT 123.190 87.520 123.360 88.220 ;
        RECT 125.330 87.520 125.500 88.220 ;
        RECT 123.575 87.290 125.115 87.460 ;
        RECT 123.190 86.530 123.360 87.230 ;
        RECT 125.330 86.530 125.500 87.230 ;
        RECT 123.575 86.300 125.115 86.470 ;
        RECT 123.190 85.540 123.360 86.240 ;
        RECT 125.330 85.540 125.500 86.240 ;
        RECT 123.575 85.310 125.115 85.480 ;
        RECT 123.190 84.550 123.360 85.250 ;
        RECT 125.330 84.550 125.500 85.250 ;
        RECT 123.575 84.320 125.115 84.490 ;
        RECT 123.190 83.560 123.360 84.260 ;
        RECT 125.330 83.560 125.500 84.260 ;
        RECT 123.575 83.330 125.115 83.500 ;
        RECT 123.190 82.570 123.360 83.270 ;
        RECT 125.330 82.570 125.500 83.270 ;
        RECT 123.575 82.340 125.115 82.510 ;
        RECT 125.840 82.200 126.250 100.470 ;
        RECT 125.840 81.940 126.010 82.200 ;
        RECT 122.680 81.770 126.010 81.940 ;
        RECT 130.510 81.940 130.680 100.730 ;
        RECT 133.670 100.330 133.840 100.730 ;
        RECT 131.405 100.160 132.945 100.330 ;
        RECT 131.020 99.400 131.190 100.100 ;
        RECT 133.160 99.400 133.330 100.100 ;
        RECT 131.405 99.170 132.945 99.340 ;
        RECT 131.020 98.410 131.190 99.110 ;
        RECT 133.160 98.410 133.330 99.110 ;
        RECT 131.405 98.180 132.945 98.350 ;
        RECT 131.020 97.420 131.190 98.120 ;
        RECT 133.160 97.420 133.330 98.120 ;
        RECT 131.405 97.190 132.945 97.360 ;
        RECT 131.020 96.430 131.190 97.130 ;
        RECT 133.160 96.430 133.330 97.130 ;
        RECT 131.405 96.200 132.945 96.370 ;
        RECT 131.020 95.440 131.190 96.140 ;
        RECT 133.160 95.440 133.330 96.140 ;
        RECT 131.405 95.210 132.945 95.380 ;
        RECT 131.020 94.450 131.190 95.150 ;
        RECT 133.160 94.450 133.330 95.150 ;
        RECT 131.405 94.220 132.945 94.390 ;
        RECT 131.020 93.460 131.190 94.160 ;
        RECT 133.160 93.460 133.330 94.160 ;
        RECT 131.405 93.230 132.945 93.400 ;
        RECT 131.020 92.470 131.190 93.170 ;
        RECT 133.160 92.470 133.330 93.170 ;
        RECT 131.405 92.240 132.945 92.410 ;
        RECT 131.020 91.480 131.190 92.180 ;
        RECT 133.160 91.480 133.330 92.180 ;
        RECT 131.405 91.250 132.945 91.420 ;
        RECT 131.020 90.490 131.190 91.190 ;
        RECT 133.160 90.490 133.330 91.190 ;
        RECT 131.405 90.260 132.945 90.430 ;
        RECT 131.020 89.500 131.190 90.200 ;
        RECT 133.160 89.500 133.330 90.200 ;
        RECT 131.405 89.270 132.945 89.440 ;
        RECT 131.020 88.510 131.190 89.210 ;
        RECT 133.160 88.510 133.330 89.210 ;
        RECT 131.405 88.280 132.945 88.450 ;
        RECT 131.020 87.520 131.190 88.220 ;
        RECT 133.160 87.520 133.330 88.220 ;
        RECT 131.405 87.290 132.945 87.460 ;
        RECT 131.020 86.530 131.190 87.230 ;
        RECT 133.160 86.530 133.330 87.230 ;
        RECT 131.405 86.300 132.945 86.470 ;
        RECT 131.020 85.540 131.190 86.240 ;
        RECT 133.160 85.540 133.330 86.240 ;
        RECT 131.405 85.310 132.945 85.480 ;
        RECT 131.020 84.550 131.190 85.250 ;
        RECT 133.160 84.550 133.330 85.250 ;
        RECT 131.405 84.320 132.945 84.490 ;
        RECT 131.020 83.560 131.190 84.260 ;
        RECT 133.160 83.560 133.330 84.260 ;
        RECT 131.405 83.330 132.945 83.500 ;
        RECT 131.020 82.570 131.190 83.270 ;
        RECT 133.160 82.570 133.330 83.270 ;
        RECT 131.405 82.340 132.945 82.510 ;
        RECT 133.660 82.230 133.960 100.330 ;
        RECT 138.350 97.360 142.180 97.530 ;
        RECT 133.670 81.940 133.840 82.230 ;
        RECT 130.510 81.770 133.840 81.940 ;
        RECT 111.910 77.770 117.650 77.940 ;
        RECT 128.040 74.140 132.010 74.310 ;
        RECT 114.900 73.630 117.640 73.800 ;
        RECT 114.900 73.360 115.070 73.630 ;
        RECT 114.840 69.060 115.070 73.360 ;
        RECT 115.750 73.060 116.790 73.230 ;
        RECT 115.410 72.000 115.580 73.000 ;
        RECT 116.960 72.000 117.130 73.000 ;
        RECT 115.750 71.770 116.790 71.940 ;
        RECT 115.410 70.710 115.580 71.710 ;
        RECT 116.960 70.710 117.130 71.710 ;
        RECT 115.750 70.480 116.790 70.650 ;
        RECT 115.410 69.420 115.580 70.420 ;
        RECT 116.960 69.420 117.130 70.420 ;
        RECT 115.750 69.190 116.790 69.360 ;
        RECT 114.900 68.790 115.070 69.060 ;
        RECT 117.470 68.790 117.640 73.630 ;
        RECT 114.900 68.620 117.640 68.790 ;
        RECT 128.040 68.690 128.210 74.140 ;
        RECT 131.840 73.890 132.010 74.140 ;
        RECT 128.935 73.570 131.115 73.740 ;
        RECT 128.550 73.160 128.720 73.510 ;
        RECT 131.330 73.160 131.500 73.510 ;
        RECT 128.935 72.930 131.115 73.100 ;
        RECT 128.550 72.520 128.720 72.870 ;
        RECT 131.330 72.520 131.500 72.870 ;
        RECT 128.935 72.290 131.115 72.460 ;
        RECT 128.550 71.880 128.720 72.230 ;
        RECT 131.330 71.880 131.500 72.230 ;
        RECT 128.935 71.650 131.115 71.820 ;
        RECT 128.550 71.240 128.720 71.590 ;
        RECT 131.330 71.240 131.500 71.590 ;
        RECT 128.935 71.010 131.115 71.180 ;
        RECT 128.550 70.600 128.720 70.950 ;
        RECT 131.330 70.600 131.500 70.950 ;
        RECT 128.935 70.370 131.115 70.540 ;
        RECT 128.550 69.960 128.720 70.310 ;
        RECT 131.330 69.960 131.500 70.310 ;
        RECT 128.935 69.730 131.115 69.900 ;
        RECT 128.550 69.320 128.720 69.670 ;
        RECT 131.330 69.320 131.500 69.670 ;
        RECT 128.935 69.090 131.115 69.260 ;
        RECT 131.840 68.940 132.100 73.890 ;
        RECT 131.840 68.690 132.010 68.940 ;
        RECT 128.040 68.520 132.010 68.690 ;
        RECT 138.350 66.780 138.520 97.360 ;
        RECT 142.010 97.080 142.180 97.360 ;
        RECT 139.245 96.790 141.285 96.960 ;
        RECT 138.860 93.730 139.030 96.730 ;
        RECT 141.500 93.730 141.670 96.730 ;
        RECT 139.245 93.500 141.285 93.670 ;
        RECT 138.860 90.440 139.030 93.440 ;
        RECT 141.500 90.440 141.670 93.440 ;
        RECT 139.245 90.210 141.285 90.380 ;
        RECT 138.860 87.150 139.030 90.150 ;
        RECT 141.500 87.150 141.670 90.150 ;
        RECT 139.245 86.920 141.285 87.090 ;
        RECT 138.860 83.860 139.030 86.860 ;
        RECT 141.500 83.860 141.670 86.860 ;
        RECT 139.245 83.630 141.285 83.800 ;
        RECT 138.860 80.570 139.030 83.570 ;
        RECT 141.500 80.570 141.670 83.570 ;
        RECT 139.245 80.340 141.285 80.510 ;
        RECT 138.860 77.280 139.030 80.280 ;
        RECT 141.500 77.280 141.670 80.280 ;
        RECT 139.245 77.050 141.285 77.220 ;
        RECT 138.860 73.990 139.030 76.990 ;
        RECT 141.500 73.990 141.670 76.990 ;
        RECT 139.245 73.760 141.285 73.930 ;
        RECT 138.860 70.700 139.030 73.700 ;
        RECT 141.500 70.700 141.670 73.700 ;
        RECT 139.245 70.470 141.285 70.640 ;
        RECT 138.860 67.410 139.030 70.410 ;
        RECT 141.500 67.410 141.670 70.410 ;
        RECT 139.245 67.180 141.285 67.350 ;
        RECT 142.010 67.040 142.250 97.080 ;
        RECT 142.010 66.780 142.180 67.040 ;
        RECT 138.350 66.610 142.180 66.780 ;
        RECT 129.170 61.110 131.910 61.280 ;
        RECT 129.170 60.860 129.340 61.110 ;
        RECT 114.930 59.660 117.670 59.830 ;
        RECT 114.930 59.410 115.100 59.660 ;
        RECT 114.780 55.070 115.100 59.410 ;
        RECT 115.780 59.090 116.820 59.260 ;
        RECT 115.440 58.030 115.610 59.030 ;
        RECT 116.990 58.030 117.160 59.030 ;
        RECT 115.780 57.800 116.820 57.970 ;
        RECT 115.440 56.740 115.610 57.740 ;
        RECT 116.990 56.740 117.160 57.740 ;
        RECT 115.780 56.510 116.820 56.680 ;
        RECT 115.440 55.450 115.610 56.450 ;
        RECT 116.990 55.450 117.160 56.450 ;
        RECT 115.780 55.220 116.820 55.390 ;
        RECT 114.930 54.820 115.100 55.070 ;
        RECT 117.500 54.820 117.670 59.660 ;
        RECT 114.930 54.650 117.670 54.820 ;
        RECT 129.100 53.500 129.340 60.860 ;
        RECT 130.020 60.540 131.060 60.710 ;
        RECT 129.680 58.480 129.850 60.480 ;
        RECT 131.230 58.480 131.400 60.480 ;
        RECT 130.020 58.250 131.060 58.420 ;
        RECT 129.680 56.190 129.850 58.190 ;
        RECT 131.230 56.190 131.400 58.190 ;
        RECT 130.020 55.960 131.060 56.130 ;
        RECT 129.680 53.900 129.850 55.900 ;
        RECT 131.230 53.900 131.400 55.900 ;
        RECT 130.020 53.670 131.060 53.840 ;
        RECT 129.170 53.270 129.340 53.500 ;
        RECT 131.740 53.270 131.910 61.110 ;
        RECT 138.000 60.280 141.500 60.450 ;
        RECT 138.000 57.390 138.170 60.280 ;
        RECT 141.330 60.020 141.500 60.280 ;
        RECT 138.895 59.710 140.605 59.880 ;
        RECT 138.510 59.300 138.680 59.650 ;
        RECT 140.820 59.300 140.990 59.650 ;
        RECT 138.895 59.070 140.605 59.240 ;
        RECT 138.510 58.660 138.680 59.010 ;
        RECT 140.820 58.660 140.990 59.010 ;
        RECT 138.895 58.430 140.605 58.600 ;
        RECT 138.510 58.020 138.680 58.370 ;
        RECT 140.820 58.020 140.990 58.370 ;
        RECT 138.895 57.790 140.605 57.960 ;
        RECT 141.330 57.650 141.580 60.020 ;
        RECT 141.330 57.390 141.500 57.650 ;
        RECT 138.000 57.220 141.500 57.390 ;
        RECT 129.170 53.100 131.910 53.270 ;
        RECT 137.800 51.720 141.630 51.890 ;
        RECT 120.700 46.240 123.440 46.410 ;
        RECT 120.700 46.010 120.870 46.240 ;
        RECT 120.470 45.060 120.870 46.010 ;
        RECT 121.210 45.370 121.380 45.700 ;
        RECT 121.550 45.670 122.590 45.840 ;
        RECT 121.550 45.230 122.590 45.400 ;
        RECT 122.760 45.370 122.930 45.700 ;
        RECT 120.700 44.830 120.870 45.060 ;
        RECT 123.270 44.830 123.440 46.240 ;
        RECT 120.700 44.660 123.440 44.830 ;
        RECT 126.030 46.290 129.860 46.460 ;
        RECT 126.030 44.680 126.200 46.290 ;
        RECT 129.690 46.050 129.860 46.290 ;
        RECT 126.925 45.720 128.965 45.890 ;
        RECT 126.540 45.310 126.710 45.660 ;
        RECT 129.180 45.310 129.350 45.660 ;
        RECT 126.925 45.080 128.965 45.250 ;
        RECT 129.690 44.940 129.960 46.050 ;
        RECT 129.690 44.680 129.860 44.940 ;
        RECT 126.030 44.510 129.860 44.680 ;
        RECT 126.030 42.150 129.860 42.320 ;
        RECT 120.700 41.560 123.940 41.730 ;
        RECT 120.700 41.320 120.870 41.560 ;
        RECT 120.450 39.870 120.870 41.320 ;
        RECT 121.210 40.670 121.380 41.000 ;
        RECT 121.550 40.990 123.090 41.160 ;
        RECT 121.550 40.510 123.090 40.680 ;
        RECT 121.550 40.030 123.090 40.200 ;
        RECT 123.260 40.190 123.430 40.520 ;
        RECT 120.700 39.630 120.870 39.870 ;
        RECT 123.770 39.630 123.940 41.560 ;
        RECT 120.700 39.460 123.940 39.630 ;
        RECT 126.030 39.260 126.200 42.150 ;
        RECT 129.690 41.900 129.860 42.150 ;
        RECT 126.925 41.580 128.965 41.750 ;
        RECT 126.540 41.170 126.710 41.520 ;
        RECT 129.180 41.170 129.350 41.520 ;
        RECT 126.925 40.940 128.965 41.110 ;
        RECT 126.540 40.530 126.710 40.880 ;
        RECT 129.180 40.530 129.350 40.880 ;
        RECT 126.925 40.300 128.965 40.470 ;
        RECT 126.540 39.890 126.710 40.240 ;
        RECT 129.180 39.890 129.350 40.240 ;
        RECT 126.925 39.660 128.965 39.830 ;
        RECT 129.690 39.500 129.930 41.900 ;
        RECT 129.690 39.260 129.860 39.500 ;
        RECT 126.030 39.090 129.860 39.260 ;
        RECT 126.030 35.930 130.860 36.100 ;
        RECT 119.260 34.730 124.000 34.900 ;
        RECT 119.260 34.470 119.430 34.730 ;
        RECT 118.940 32.570 119.430 34.470 ;
        RECT 119.770 33.840 119.940 34.170 ;
        RECT 120.110 34.160 123.150 34.330 ;
        RECT 120.110 33.680 123.150 33.850 ;
        RECT 119.770 32.880 119.940 33.210 ;
        RECT 120.110 33.200 123.150 33.370 ;
        RECT 123.320 33.360 123.490 33.690 ;
        RECT 120.110 32.720 123.150 32.890 ;
        RECT 119.260 32.320 119.430 32.570 ;
        RECT 123.830 32.320 124.000 34.730 ;
        RECT 119.260 32.150 124.000 32.320 ;
        RECT 126.030 31.120 126.200 35.930 ;
        RECT 130.690 35.670 130.860 35.930 ;
        RECT 126.925 35.360 129.965 35.530 ;
        RECT 126.540 34.950 126.710 35.300 ;
        RECT 130.180 34.950 130.350 35.300 ;
        RECT 126.925 34.720 129.965 34.890 ;
        RECT 126.540 34.310 126.710 34.660 ;
        RECT 130.180 34.310 130.350 34.660 ;
        RECT 126.925 34.080 129.965 34.250 ;
        RECT 126.540 33.670 126.710 34.020 ;
        RECT 130.180 33.670 130.350 34.020 ;
        RECT 126.925 33.440 129.965 33.610 ;
        RECT 126.540 33.030 126.710 33.380 ;
        RECT 130.180 33.030 130.350 33.380 ;
        RECT 126.925 32.800 129.965 32.970 ;
        RECT 126.540 32.390 126.710 32.740 ;
        RECT 130.180 32.390 130.350 32.740 ;
        RECT 126.925 32.160 129.965 32.330 ;
        RECT 126.540 31.750 126.710 32.100 ;
        RECT 130.180 31.750 130.350 32.100 ;
        RECT 126.925 31.520 129.965 31.690 ;
        RECT 130.690 31.390 130.920 35.670 ;
        RECT 130.690 31.120 130.860 31.390 ;
        RECT 126.030 30.950 130.860 31.120 ;
        RECT 137.800 31.010 137.970 51.720 ;
        RECT 141.460 51.450 141.630 51.720 ;
        RECT 138.695 51.150 140.735 51.320 ;
        RECT 138.310 48.090 138.480 51.090 ;
        RECT 140.950 48.090 141.120 51.090 ;
        RECT 138.695 47.860 140.735 48.030 ;
        RECT 138.310 44.800 138.480 47.800 ;
        RECT 140.950 44.800 141.120 47.800 ;
        RECT 138.695 44.570 140.735 44.740 ;
        RECT 138.310 41.510 138.480 44.510 ;
        RECT 140.950 41.510 141.120 44.510 ;
        RECT 138.695 41.280 140.735 41.450 ;
        RECT 138.310 38.220 138.480 41.220 ;
        RECT 140.950 38.220 141.120 41.220 ;
        RECT 138.695 37.990 140.735 38.160 ;
        RECT 138.310 34.930 138.480 37.930 ;
        RECT 140.950 34.930 141.120 37.930 ;
        RECT 138.695 34.700 140.735 34.870 ;
        RECT 138.310 31.640 138.480 34.640 ;
        RECT 140.950 31.640 141.120 34.640 ;
        RECT 138.695 31.410 140.735 31.580 ;
        RECT 141.460 31.270 141.710 51.450 ;
        RECT 141.460 31.010 141.630 31.270 ;
        RECT 137.800 30.840 141.630 31.010 ;
      LAYER mcon ;
        RECT 112.200 118.980 115.080 119.150 ;
        RECT 111.780 116.000 111.950 118.840 ;
        RECT 115.330 116.000 115.500 118.840 ;
        RECT 112.200 115.690 115.080 115.860 ;
        RECT 121.380 119.550 125.230 119.770 ;
        RECT 121.860 118.980 124.740 119.150 ;
        RECT 121.440 118.740 121.610 118.910 ;
        RECT 121.860 118.500 124.740 118.670 ;
        RECT 124.990 118.260 125.160 118.430 ;
        RECT 121.860 118.020 124.740 118.190 ;
        RECT 121.440 117.780 121.610 117.950 ;
        RECT 121.860 117.540 124.740 117.710 ;
        RECT 124.990 117.300 125.160 117.470 ;
        RECT 121.860 117.060 124.740 117.230 ;
        RECT 121.440 116.820 121.610 116.990 ;
        RECT 121.860 116.580 124.740 116.750 ;
        RECT 124.990 116.340 125.160 116.510 ;
        RECT 121.860 116.100 124.740 116.270 ;
        RECT 121.440 115.860 121.610 116.030 ;
        RECT 121.860 115.620 124.740 115.790 ;
        RECT 130.520 119.550 134.420 119.750 ;
        RECT 131.035 118.980 133.915 119.150 ;
        RECT 130.570 118.650 130.740 118.840 ;
        RECT 134.210 118.650 134.380 118.840 ;
        RECT 131.035 118.340 133.915 118.510 ;
        RECT 130.570 118.010 130.740 118.200 ;
        RECT 134.210 118.010 134.380 118.200 ;
        RECT 131.035 117.700 133.915 117.870 ;
        RECT 130.570 117.370 130.740 117.560 ;
        RECT 134.210 117.370 134.380 117.560 ;
        RECT 131.035 117.060 133.915 117.230 ;
        RECT 130.570 116.730 130.740 116.920 ;
        RECT 134.210 116.730 134.380 116.920 ;
        RECT 131.035 116.420 133.915 116.590 ;
        RECT 130.570 116.090 130.740 116.280 ;
        RECT 134.210 116.090 134.380 116.280 ;
        RECT 131.035 115.780 133.915 115.950 ;
        RECT 130.570 115.450 130.740 115.640 ;
        RECT 134.210 115.450 134.380 115.640 ;
        RECT 131.035 115.140 133.915 115.310 ;
        RECT 130.570 114.810 130.740 115.000 ;
        RECT 134.210 114.810 134.380 115.000 ;
        RECT 131.035 114.500 133.915 114.670 ;
        RECT 139.425 118.870 142.305 119.040 ;
        RECT 138.960 115.890 139.130 118.730 ;
        RECT 142.600 115.890 142.770 118.730 ;
        RECT 139.425 115.580 142.305 115.750 ;
        RECT 112.780 103.810 116.660 103.980 ;
        RECT 112.360 100.830 112.530 103.670 ;
        RECT 116.910 100.830 117.080 103.670 ;
        RECT 112.780 100.520 116.660 100.690 ;
        RECT 112.360 97.540 112.530 100.380 ;
        RECT 116.910 97.540 117.080 100.380 ;
        RECT 112.780 97.230 116.660 97.400 ;
        RECT 112.360 94.250 112.530 97.090 ;
        RECT 116.910 94.250 117.080 97.090 ;
        RECT 112.780 93.940 116.660 94.110 ;
        RECT 112.840 88.210 116.720 88.380 ;
        RECT 112.420 85.230 112.590 88.070 ;
        RECT 116.970 85.230 117.140 88.070 ;
        RECT 112.840 84.920 116.720 85.090 ;
        RECT 112.420 81.940 112.590 84.780 ;
        RECT 116.970 81.940 117.140 84.780 ;
        RECT 112.840 81.630 116.720 81.800 ;
        RECT 112.420 78.650 112.590 81.490 ;
        RECT 116.970 78.650 117.140 81.490 ;
        RECT 112.840 78.340 116.720 78.510 ;
        RECT 123.655 100.160 125.035 100.330 ;
        RECT 123.190 99.480 123.360 100.020 ;
        RECT 125.330 99.480 125.500 100.020 ;
        RECT 123.655 99.170 125.035 99.340 ;
        RECT 123.190 98.490 123.360 99.030 ;
        RECT 125.330 98.490 125.500 99.030 ;
        RECT 123.655 98.180 125.035 98.350 ;
        RECT 123.190 97.500 123.360 98.040 ;
        RECT 125.330 97.500 125.500 98.040 ;
        RECT 123.655 97.190 125.035 97.360 ;
        RECT 123.190 96.510 123.360 97.050 ;
        RECT 125.330 96.510 125.500 97.050 ;
        RECT 123.655 96.200 125.035 96.370 ;
        RECT 123.190 95.520 123.360 96.060 ;
        RECT 125.330 95.520 125.500 96.060 ;
        RECT 123.655 95.210 125.035 95.380 ;
        RECT 123.190 94.530 123.360 95.070 ;
        RECT 125.330 94.530 125.500 95.070 ;
        RECT 123.655 94.220 125.035 94.390 ;
        RECT 123.190 93.540 123.360 94.080 ;
        RECT 125.330 93.540 125.500 94.080 ;
        RECT 123.655 93.230 125.035 93.400 ;
        RECT 123.190 92.550 123.360 93.090 ;
        RECT 125.330 92.550 125.500 93.090 ;
        RECT 123.655 92.240 125.035 92.410 ;
        RECT 123.190 91.560 123.360 92.100 ;
        RECT 125.330 91.560 125.500 92.100 ;
        RECT 123.655 91.250 125.035 91.420 ;
        RECT 123.190 90.570 123.360 91.110 ;
        RECT 125.330 90.570 125.500 91.110 ;
        RECT 123.655 90.260 125.035 90.430 ;
        RECT 123.190 89.580 123.360 90.120 ;
        RECT 125.330 89.580 125.500 90.120 ;
        RECT 123.655 89.270 125.035 89.440 ;
        RECT 123.190 88.590 123.360 89.130 ;
        RECT 125.330 88.590 125.500 89.130 ;
        RECT 123.655 88.280 125.035 88.450 ;
        RECT 123.190 87.600 123.360 88.140 ;
        RECT 125.330 87.600 125.500 88.140 ;
        RECT 123.655 87.290 125.035 87.460 ;
        RECT 123.190 86.610 123.360 87.150 ;
        RECT 125.330 86.610 125.500 87.150 ;
        RECT 123.655 86.300 125.035 86.470 ;
        RECT 123.190 85.620 123.360 86.160 ;
        RECT 125.330 85.620 125.500 86.160 ;
        RECT 123.655 85.310 125.035 85.480 ;
        RECT 123.190 84.630 123.360 85.170 ;
        RECT 125.330 84.630 125.500 85.170 ;
        RECT 123.655 84.320 125.035 84.490 ;
        RECT 123.190 83.640 123.360 84.180 ;
        RECT 125.330 83.640 125.500 84.180 ;
        RECT 123.655 83.330 125.035 83.500 ;
        RECT 123.190 82.650 123.360 83.190 ;
        RECT 125.330 82.650 125.500 83.190 ;
        RECT 123.655 82.340 125.035 82.510 ;
        RECT 131.485 100.160 132.865 100.330 ;
        RECT 131.020 99.480 131.190 100.020 ;
        RECT 133.160 99.480 133.330 100.020 ;
        RECT 131.485 99.170 132.865 99.340 ;
        RECT 131.020 98.490 131.190 99.030 ;
        RECT 133.160 98.490 133.330 99.030 ;
        RECT 131.485 98.180 132.865 98.350 ;
        RECT 131.020 97.500 131.190 98.040 ;
        RECT 133.160 97.500 133.330 98.040 ;
        RECT 131.485 97.190 132.865 97.360 ;
        RECT 131.020 96.510 131.190 97.050 ;
        RECT 133.160 96.510 133.330 97.050 ;
        RECT 131.485 96.200 132.865 96.370 ;
        RECT 131.020 95.520 131.190 96.060 ;
        RECT 133.160 95.520 133.330 96.060 ;
        RECT 131.485 95.210 132.865 95.380 ;
        RECT 131.020 94.530 131.190 95.070 ;
        RECT 133.160 94.530 133.330 95.070 ;
        RECT 131.485 94.220 132.865 94.390 ;
        RECT 131.020 93.540 131.190 94.080 ;
        RECT 133.160 93.540 133.330 94.080 ;
        RECT 131.485 93.230 132.865 93.400 ;
        RECT 131.020 92.550 131.190 93.090 ;
        RECT 133.160 92.550 133.330 93.090 ;
        RECT 131.485 92.240 132.865 92.410 ;
        RECT 131.020 91.560 131.190 92.100 ;
        RECT 133.160 91.560 133.330 92.100 ;
        RECT 131.485 91.250 132.865 91.420 ;
        RECT 131.020 90.570 131.190 91.110 ;
        RECT 133.160 90.570 133.330 91.110 ;
        RECT 131.485 90.260 132.865 90.430 ;
        RECT 131.020 89.580 131.190 90.120 ;
        RECT 133.160 89.580 133.330 90.120 ;
        RECT 131.485 89.270 132.865 89.440 ;
        RECT 131.020 88.590 131.190 89.130 ;
        RECT 133.160 88.590 133.330 89.130 ;
        RECT 131.485 88.280 132.865 88.450 ;
        RECT 131.020 87.600 131.190 88.140 ;
        RECT 133.160 87.600 133.330 88.140 ;
        RECT 131.485 87.290 132.865 87.460 ;
        RECT 131.020 86.610 131.190 87.150 ;
        RECT 133.160 86.610 133.330 87.150 ;
        RECT 131.485 86.300 132.865 86.470 ;
        RECT 131.020 85.620 131.190 86.160 ;
        RECT 133.160 85.620 133.330 86.160 ;
        RECT 131.485 85.310 132.865 85.480 ;
        RECT 131.020 84.630 131.190 85.170 ;
        RECT 133.160 84.630 133.330 85.170 ;
        RECT 131.485 84.320 132.865 84.490 ;
        RECT 131.020 83.640 131.190 84.180 ;
        RECT 133.160 83.640 133.330 84.180 ;
        RECT 131.485 83.330 132.865 83.500 ;
        RECT 131.020 82.650 131.190 83.190 ;
        RECT 133.160 82.650 133.330 83.190 ;
        RECT 131.485 82.340 132.865 82.510 ;
        RECT 115.830 73.060 116.710 73.230 ;
        RECT 115.410 72.080 115.580 72.920 ;
        RECT 116.960 72.080 117.130 72.920 ;
        RECT 115.830 71.770 116.710 71.940 ;
        RECT 115.410 70.790 115.580 71.630 ;
        RECT 116.960 70.790 117.130 71.630 ;
        RECT 115.830 70.480 116.710 70.650 ;
        RECT 115.410 69.500 115.580 70.340 ;
        RECT 116.960 69.500 117.130 70.340 ;
        RECT 115.830 69.190 116.710 69.360 ;
        RECT 129.015 73.570 131.035 73.740 ;
        RECT 128.550 73.240 128.720 73.430 ;
        RECT 131.330 73.240 131.500 73.430 ;
        RECT 129.015 72.930 131.035 73.100 ;
        RECT 128.550 72.600 128.720 72.790 ;
        RECT 131.330 72.600 131.500 72.790 ;
        RECT 129.015 72.290 131.035 72.460 ;
        RECT 128.550 71.960 128.720 72.150 ;
        RECT 131.330 71.960 131.500 72.150 ;
        RECT 129.015 71.650 131.035 71.820 ;
        RECT 128.550 71.320 128.720 71.510 ;
        RECT 131.330 71.320 131.500 71.510 ;
        RECT 129.015 71.010 131.035 71.180 ;
        RECT 128.550 70.680 128.720 70.870 ;
        RECT 131.330 70.680 131.500 70.870 ;
        RECT 129.015 70.370 131.035 70.540 ;
        RECT 128.550 70.040 128.720 70.230 ;
        RECT 131.330 70.040 131.500 70.230 ;
        RECT 129.015 69.730 131.035 69.900 ;
        RECT 128.550 69.400 128.720 69.590 ;
        RECT 131.330 69.400 131.500 69.590 ;
        RECT 129.015 69.090 131.035 69.260 ;
        RECT 139.325 96.790 141.205 96.960 ;
        RECT 138.860 93.810 139.030 96.650 ;
        RECT 141.500 93.810 141.670 96.650 ;
        RECT 139.325 93.500 141.205 93.670 ;
        RECT 138.860 90.520 139.030 93.360 ;
        RECT 141.500 90.520 141.670 93.360 ;
        RECT 139.325 90.210 141.205 90.380 ;
        RECT 138.860 87.230 139.030 90.070 ;
        RECT 141.500 87.230 141.670 90.070 ;
        RECT 139.325 86.920 141.205 87.090 ;
        RECT 138.860 83.940 139.030 86.780 ;
        RECT 141.500 83.940 141.670 86.780 ;
        RECT 139.325 83.630 141.205 83.800 ;
        RECT 138.860 80.650 139.030 83.490 ;
        RECT 141.500 80.650 141.670 83.490 ;
        RECT 139.325 80.340 141.205 80.510 ;
        RECT 138.860 77.360 139.030 80.200 ;
        RECT 141.500 77.360 141.670 80.200 ;
        RECT 139.325 77.050 141.205 77.220 ;
        RECT 138.860 74.070 139.030 76.910 ;
        RECT 141.500 74.070 141.670 76.910 ;
        RECT 139.325 73.760 141.205 73.930 ;
        RECT 138.860 70.780 139.030 73.620 ;
        RECT 141.500 70.780 141.670 73.620 ;
        RECT 139.325 70.470 141.205 70.640 ;
        RECT 138.860 67.490 139.030 70.330 ;
        RECT 141.500 67.490 141.670 70.330 ;
        RECT 139.325 67.180 141.205 67.350 ;
        RECT 115.860 59.090 116.740 59.260 ;
        RECT 115.440 58.110 115.610 58.950 ;
        RECT 116.990 58.110 117.160 58.950 ;
        RECT 115.860 57.800 116.740 57.970 ;
        RECT 115.440 56.820 115.610 57.660 ;
        RECT 116.990 56.820 117.160 57.660 ;
        RECT 115.860 56.510 116.740 56.680 ;
        RECT 115.440 55.530 115.610 56.370 ;
        RECT 116.990 55.530 117.160 56.370 ;
        RECT 115.860 55.220 116.740 55.390 ;
        RECT 130.100 60.540 130.980 60.710 ;
        RECT 129.680 58.560 129.850 60.400 ;
        RECT 131.230 58.560 131.400 60.400 ;
        RECT 130.100 58.250 130.980 58.420 ;
        RECT 129.680 56.270 129.850 58.110 ;
        RECT 131.230 56.270 131.400 58.110 ;
        RECT 130.100 55.960 130.980 56.130 ;
        RECT 129.680 53.980 129.850 55.820 ;
        RECT 131.230 53.980 131.400 55.820 ;
        RECT 130.100 53.670 130.980 53.840 ;
        RECT 138.975 59.710 140.525 59.880 ;
        RECT 138.510 59.380 138.680 59.570 ;
        RECT 140.820 59.380 140.990 59.570 ;
        RECT 138.975 59.070 140.525 59.240 ;
        RECT 138.510 58.740 138.680 58.930 ;
        RECT 140.820 58.740 140.990 58.930 ;
        RECT 138.975 58.430 140.525 58.600 ;
        RECT 138.510 58.100 138.680 58.290 ;
        RECT 140.820 58.100 140.990 58.290 ;
        RECT 138.975 57.790 140.525 57.960 ;
        RECT 121.630 45.670 122.510 45.840 ;
        RECT 121.210 45.450 121.380 45.620 ;
        RECT 122.760 45.450 122.930 45.620 ;
        RECT 121.630 45.230 122.510 45.400 ;
        RECT 127.005 45.720 128.885 45.890 ;
        RECT 126.540 45.390 126.710 45.580 ;
        RECT 129.180 45.390 129.350 45.580 ;
        RECT 127.005 45.080 128.885 45.250 ;
        RECT 121.630 40.990 123.010 41.160 ;
        RECT 121.210 40.750 121.380 40.920 ;
        RECT 121.630 40.510 123.010 40.680 ;
        RECT 123.260 40.270 123.430 40.440 ;
        RECT 121.630 40.030 123.010 40.200 ;
        RECT 127.005 41.580 128.885 41.750 ;
        RECT 126.540 41.250 126.710 41.440 ;
        RECT 129.180 41.250 129.350 41.440 ;
        RECT 127.005 40.940 128.885 41.110 ;
        RECT 126.540 40.610 126.710 40.800 ;
        RECT 129.180 40.610 129.350 40.800 ;
        RECT 127.005 40.300 128.885 40.470 ;
        RECT 126.540 39.970 126.710 40.160 ;
        RECT 129.180 39.970 129.350 40.160 ;
        RECT 127.005 39.660 128.885 39.830 ;
        RECT 120.190 34.160 123.070 34.330 ;
        RECT 119.770 33.920 119.940 34.090 ;
        RECT 120.190 33.680 123.070 33.850 ;
        RECT 123.320 33.440 123.490 33.610 ;
        RECT 120.190 33.200 123.070 33.370 ;
        RECT 119.770 32.960 119.940 33.130 ;
        RECT 120.190 32.720 123.070 32.890 ;
        RECT 127.005 35.360 129.885 35.530 ;
        RECT 126.540 35.030 126.710 35.220 ;
        RECT 130.180 35.030 130.350 35.220 ;
        RECT 127.005 34.720 129.885 34.890 ;
        RECT 126.540 34.390 126.710 34.580 ;
        RECT 130.180 34.390 130.350 34.580 ;
        RECT 127.005 34.080 129.885 34.250 ;
        RECT 126.540 33.750 126.710 33.940 ;
        RECT 130.180 33.750 130.350 33.940 ;
        RECT 127.005 33.440 129.885 33.610 ;
        RECT 126.540 33.110 126.710 33.300 ;
        RECT 130.180 33.110 130.350 33.300 ;
        RECT 127.005 32.800 129.885 32.970 ;
        RECT 126.540 32.470 126.710 32.660 ;
        RECT 130.180 32.470 130.350 32.660 ;
        RECT 127.005 32.160 129.885 32.330 ;
        RECT 126.540 31.830 126.710 32.020 ;
        RECT 130.180 31.830 130.350 32.020 ;
        RECT 127.005 31.520 129.885 31.690 ;
        RECT 138.775 51.150 140.655 51.320 ;
        RECT 138.310 48.170 138.480 51.010 ;
        RECT 140.950 48.170 141.120 51.010 ;
        RECT 138.775 47.860 140.655 48.030 ;
        RECT 138.310 44.880 138.480 47.720 ;
        RECT 140.950 44.880 141.120 47.720 ;
        RECT 138.775 44.570 140.655 44.740 ;
        RECT 138.310 41.590 138.480 44.430 ;
        RECT 140.950 41.590 141.120 44.430 ;
        RECT 138.775 41.280 140.655 41.450 ;
        RECT 138.310 38.300 138.480 41.140 ;
        RECT 140.950 38.300 141.120 41.140 ;
        RECT 138.775 37.990 140.655 38.160 ;
        RECT 138.310 35.010 138.480 37.850 ;
        RECT 140.950 35.010 141.120 37.850 ;
        RECT 138.775 34.700 140.655 34.870 ;
        RECT 138.310 31.720 138.480 34.560 ;
        RECT 140.950 31.720 141.120 34.560 ;
        RECT 138.775 31.410 140.655 31.580 ;
        RECT 141.470 31.270 141.710 51.450 ;
      LAYER met1 ;
        RECT 86.900 134.210 88.400 134.240 ;
        RECT 106.900 134.225 108.680 134.350 ;
        RECT 102.965 134.210 108.680 134.225 ;
        RECT 86.900 132.710 108.680 134.210 ;
        RECT 86.900 132.680 88.400 132.710 ;
        RECT 102.965 132.695 108.680 132.710 ;
        RECT 106.900 124.300 108.680 132.695 ;
        RECT 127.360 128.760 137.935 130.025 ;
        RECT 127.360 124.650 128.625 128.760 ;
        RECT 106.010 124.290 110.030 124.300 ;
        RECT 106.010 122.010 125.510 124.290 ;
        RECT 106.010 121.930 125.520 122.010 ;
        RECT 106.010 119.530 110.030 121.930 ;
        RECT 106.010 115.290 111.470 119.530 ;
        RECT 112.180 119.180 115.110 121.930 ;
        RECT 121.190 119.520 125.520 121.930 ;
        RECT 124.310 119.180 124.800 119.240 ;
        RECT 112.140 118.950 115.140 119.180 ;
        RECT 106.010 104.160 110.030 115.290 ;
        RECT 111.750 112.730 111.990 118.920 ;
        RECT 112.210 115.890 115.110 115.910 ;
        RECT 112.140 115.660 115.140 115.890 ;
        RECT 112.210 115.490 115.110 115.660 ;
        RECT 112.860 114.660 113.700 115.490 ;
        RECT 112.865 112.730 113.695 114.660 ;
        RECT 115.290 112.730 115.590 118.930 ;
        RECT 118.940 113.940 119.560 114.500 ;
        RECT 118.970 112.730 119.530 113.940 ;
        RECT 111.750 112.130 119.530 112.730 ;
        RECT 121.290 112.690 121.640 119.000 ;
        RECT 121.800 118.950 124.800 119.180 ;
        RECT 124.310 118.850 124.800 118.950 ;
        RECT 121.870 118.700 122.360 118.780 ;
        RECT 121.800 118.470 124.800 118.700 ;
        RECT 121.870 118.390 122.360 118.470 ;
        RECT 124.310 118.220 124.800 118.300 ;
        RECT 121.800 117.990 124.800 118.220 ;
        RECT 124.310 117.910 124.800 117.990 ;
        RECT 121.870 117.740 122.360 117.820 ;
        RECT 121.800 117.510 124.800 117.740 ;
        RECT 121.870 117.430 122.360 117.510 ;
        RECT 124.310 117.260 124.800 117.340 ;
        RECT 121.800 117.030 124.800 117.260 ;
        RECT 124.310 116.950 124.800 117.030 ;
        RECT 121.870 116.780 122.360 116.860 ;
        RECT 121.800 116.550 124.800 116.780 ;
        RECT 121.870 116.470 122.360 116.550 ;
        RECT 124.310 116.300 124.800 116.380 ;
        RECT 121.800 116.070 124.800 116.300 ;
        RECT 124.310 115.990 124.800 116.070 ;
        RECT 121.870 115.820 122.360 115.900 ;
        RECT 121.800 115.590 124.800 115.820 ;
        RECT 121.870 115.510 122.360 115.590 ;
        RECT 123.495 112.690 124.065 114.590 ;
        RECT 124.940 112.690 125.290 118.550 ;
        RECT 127.230 115.400 128.795 124.650 ;
        RECT 144.960 124.440 146.825 143.225 ;
        RECT 130.450 122.150 148.100 124.440 ;
        RECT 130.440 122.080 148.100 122.150 ;
        RECT 130.440 119.480 134.460 122.080 ;
        RECT 131.050 119.180 131.530 119.190 ;
        RECT 130.470 113.310 130.780 118.980 ;
        RECT 130.975 118.950 133.975 119.180 ;
        RECT 139.560 119.070 142.090 122.080 ;
        RECT 144.080 119.610 148.100 122.080 ;
        RECT 131.050 118.810 131.530 118.950 ;
        RECT 133.450 118.540 133.930 118.620 ;
        RECT 130.975 118.310 133.975 118.540 ;
        RECT 133.450 118.240 133.930 118.310 ;
        RECT 131.030 117.900 131.510 117.970 ;
        RECT 130.975 117.670 133.975 117.900 ;
        RECT 131.030 117.590 131.510 117.670 ;
        RECT 133.450 117.260 133.930 117.330 ;
        RECT 130.975 117.030 133.975 117.260 ;
        RECT 133.450 116.950 133.930 117.030 ;
        RECT 131.030 116.620 131.510 116.700 ;
        RECT 130.975 116.390 133.975 116.620 ;
        RECT 131.030 116.320 131.510 116.390 ;
        RECT 133.450 115.980 133.930 116.060 ;
        RECT 130.975 115.750 133.975 115.980 ;
        RECT 133.450 115.680 133.930 115.750 ;
        RECT 131.030 115.340 131.510 115.410 ;
        RECT 130.975 115.110 133.975 115.340 ;
        RECT 131.030 115.030 131.510 115.110 ;
        RECT 133.450 114.700 133.930 114.780 ;
        RECT 130.975 114.470 133.975 114.700 ;
        RECT 133.450 114.400 133.930 114.470 ;
        RECT 130.470 112.730 131.610 113.310 ;
        RECT 130.470 112.690 131.580 112.730 ;
        RECT 121.280 112.420 131.580 112.690 ;
        RECT 134.130 112.420 134.440 118.980 ;
        RECT 138.890 118.790 139.140 118.870 ;
        RECT 139.365 118.840 142.365 119.070 ;
        RECT 142.540 118.790 142.790 118.870 ;
        RECT 138.890 115.830 139.160 118.790 ;
        RECT 142.540 115.830 142.800 118.790 ;
        RECT 138.890 114.180 139.140 115.830 ;
        RECT 139.365 115.550 142.365 115.780 ;
        RECT 140.510 114.180 141.660 115.550 ;
        RECT 142.540 114.180 142.790 115.830 ;
        RECT 143.080 114.990 148.100 119.610 ;
        RECT 138.890 114.005 142.790 114.180 ;
        RECT 136.795 113.455 142.795 114.005 ;
        RECT 135.920 113.270 136.460 113.300 ;
        RECT 136.795 113.270 137.345 113.455 ;
        RECT 135.920 112.730 137.345 113.270 ;
        RECT 135.920 112.700 136.460 112.730 ;
        RECT 136.795 112.725 137.345 112.730 ;
        RECT 111.750 112.050 119.510 112.130 ;
        RECT 121.280 112.110 134.445 112.420 ;
        RECT 121.280 112.090 130.920 112.110 ;
        RECT 116.280 109.540 117.210 112.050 ;
        RECT 141.110 110.365 141.700 113.455 ;
        RECT 141.080 109.775 141.730 110.365 ;
        RECT 116.280 108.600 120.210 109.540 ;
        RECT 116.280 107.530 117.210 108.600 ;
        RECT 112.330 106.090 117.220 107.530 ;
        RECT 106.010 93.720 112.050 104.160 ;
        RECT 112.330 94.160 112.580 106.090 ;
        RECT 116.020 104.010 116.650 104.100 ;
        RECT 112.720 103.780 116.720 104.010 ;
        RECT 116.020 103.680 116.650 103.780 ;
        RECT 112.790 100.720 113.420 100.830 ;
        RECT 112.720 100.490 116.720 100.720 ;
        RECT 112.790 100.410 113.420 100.490 ;
        RECT 116.020 97.430 116.650 97.520 ;
        RECT 112.720 97.200 116.720 97.430 ;
        RECT 116.020 97.100 116.650 97.200 ;
        RECT 112.790 94.140 113.420 94.220 ;
        RECT 112.720 93.910 116.720 94.140 ;
        RECT 116.880 93.960 117.220 106.090 ;
        RECT 112.790 93.800 113.420 93.910 ;
        RECT 106.010 92.540 110.030 93.720 ;
        RECT 106.010 91.790 113.520 92.540 ;
        RECT 106.010 88.710 110.030 91.790 ;
        RECT 116.930 90.430 117.310 90.440 ;
        RECT 119.270 90.430 120.210 108.600 ;
        RECT 126.250 105.480 127.640 105.485 ;
        RECT 133.960 105.480 135.550 105.485 ;
        RECT 144.080 105.480 148.100 114.990 ;
        RECT 126.250 102.260 148.100 105.480 ;
        RECT 126.250 100.580 127.640 102.260 ;
        RECT 124.630 100.360 125.040 100.440 ;
        RECT 112.390 89.490 120.210 90.430 ;
        RECT 106.010 78.110 112.110 88.710 ;
        RECT 112.390 78.590 112.640 89.490 ;
        RECT 116.020 88.410 116.730 88.520 ;
        RECT 112.780 88.180 116.780 88.410 ;
        RECT 116.020 88.050 116.730 88.180 ;
        RECT 112.840 85.120 113.550 85.230 ;
        RECT 112.780 84.890 116.780 85.120 ;
        RECT 112.840 84.760 113.550 84.890 ;
        RECT 116.020 81.830 116.730 81.950 ;
        RECT 112.780 81.600 116.780 81.830 ;
        RECT 116.020 81.480 116.730 81.600 ;
        RECT 112.840 78.540 113.550 78.660 ;
        RECT 112.780 78.310 116.780 78.540 ;
        RECT 116.930 78.470 117.310 89.490 ;
        RECT 123.090 80.670 123.410 100.160 ;
        RECT 123.595 100.130 125.095 100.360 ;
        RECT 124.630 100.050 125.040 100.130 ;
        RECT 123.650 99.370 124.060 99.450 ;
        RECT 123.595 99.140 125.095 99.370 ;
        RECT 123.650 99.060 124.060 99.140 ;
        RECT 124.630 98.380 125.040 98.460 ;
        RECT 123.595 98.150 125.095 98.380 ;
        RECT 124.630 98.070 125.040 98.150 ;
        RECT 123.650 97.390 124.060 97.470 ;
        RECT 123.595 97.160 125.095 97.390 ;
        RECT 123.650 97.080 124.060 97.160 ;
        RECT 124.630 96.400 125.040 96.480 ;
        RECT 123.595 96.170 125.095 96.400 ;
        RECT 124.630 96.090 125.040 96.170 ;
        RECT 123.650 95.410 124.060 95.490 ;
        RECT 123.595 95.180 125.095 95.410 ;
        RECT 123.650 95.100 124.060 95.180 ;
        RECT 124.630 94.420 125.040 94.500 ;
        RECT 123.595 94.190 125.095 94.420 ;
        RECT 124.630 94.110 125.040 94.190 ;
        RECT 123.650 93.430 124.060 93.520 ;
        RECT 123.595 93.200 125.095 93.430 ;
        RECT 123.650 93.130 124.060 93.200 ;
        RECT 124.630 92.440 125.040 92.520 ;
        RECT 123.595 92.210 125.095 92.440 ;
        RECT 124.630 92.130 125.040 92.210 ;
        RECT 123.650 91.450 124.060 91.540 ;
        RECT 123.595 91.220 125.095 91.450 ;
        RECT 123.650 91.150 124.060 91.220 ;
        RECT 124.630 90.460 125.040 90.540 ;
        RECT 123.595 90.230 125.095 90.460 ;
        RECT 124.630 90.150 125.040 90.230 ;
        RECT 123.650 89.470 124.060 89.550 ;
        RECT 123.595 89.240 125.095 89.470 ;
        RECT 123.650 89.160 124.060 89.240 ;
        RECT 124.630 88.480 125.040 88.560 ;
        RECT 123.595 88.250 125.095 88.480 ;
        RECT 124.630 88.170 125.040 88.250 ;
        RECT 123.650 87.490 124.060 87.580 ;
        RECT 123.595 87.260 125.095 87.490 ;
        RECT 123.650 87.190 124.060 87.260 ;
        RECT 124.630 86.500 125.040 86.580 ;
        RECT 123.595 86.270 125.095 86.500 ;
        RECT 124.630 86.190 125.040 86.270 ;
        RECT 123.650 85.510 124.060 85.590 ;
        RECT 123.595 85.280 125.095 85.510 ;
        RECT 123.650 85.200 124.060 85.280 ;
        RECT 124.630 84.520 125.040 84.600 ;
        RECT 123.595 84.290 125.095 84.520 ;
        RECT 124.630 84.210 125.040 84.290 ;
        RECT 123.650 83.530 124.060 83.610 ;
        RECT 123.595 83.300 125.095 83.530 ;
        RECT 123.650 83.220 124.060 83.300 ;
        RECT 124.630 82.540 125.040 82.620 ;
        RECT 123.595 82.310 125.095 82.540 ;
        RECT 124.630 82.230 125.040 82.310 ;
        RECT 125.250 80.670 125.570 100.160 ;
        RECT 125.780 82.030 127.640 100.580 ;
        RECT 133.960 100.460 135.550 102.260 ;
        RECT 132.420 100.360 132.950 100.440 ;
        RECT 131.425 100.130 132.950 100.360 ;
        RECT 130.910 80.670 131.230 100.100 ;
        RECT 132.420 100.050 132.950 100.130 ;
        RECT 131.460 99.370 131.990 99.450 ;
        RECT 131.425 99.140 132.925 99.370 ;
        RECT 131.460 99.060 131.990 99.140 ;
        RECT 132.420 98.380 132.950 98.460 ;
        RECT 131.425 98.150 132.950 98.380 ;
        RECT 132.420 98.070 132.950 98.150 ;
        RECT 131.460 97.390 131.990 97.480 ;
        RECT 131.425 97.160 132.925 97.390 ;
        RECT 131.460 97.090 131.990 97.160 ;
        RECT 132.420 96.400 132.950 96.480 ;
        RECT 131.425 96.170 132.950 96.400 ;
        RECT 132.420 96.090 132.950 96.170 ;
        RECT 131.460 95.410 131.990 95.500 ;
        RECT 131.425 95.180 132.925 95.410 ;
        RECT 131.460 95.110 131.990 95.180 ;
        RECT 132.420 94.420 132.950 94.510 ;
        RECT 131.425 94.190 132.950 94.420 ;
        RECT 132.420 94.120 132.950 94.190 ;
        RECT 131.460 93.430 131.990 93.510 ;
        RECT 131.425 93.200 132.925 93.430 ;
        RECT 131.460 93.120 131.990 93.200 ;
        RECT 132.420 92.440 132.950 92.530 ;
        RECT 131.425 92.210 132.950 92.440 ;
        RECT 132.420 92.140 132.950 92.210 ;
        RECT 131.460 91.450 131.990 91.530 ;
        RECT 131.425 91.220 132.925 91.450 ;
        RECT 131.460 91.140 131.990 91.220 ;
        RECT 132.420 90.460 132.950 90.540 ;
        RECT 131.425 90.230 132.950 90.460 ;
        RECT 132.420 90.150 132.950 90.230 ;
        RECT 131.460 89.470 131.990 89.560 ;
        RECT 131.425 89.240 132.925 89.470 ;
        RECT 131.460 89.170 131.990 89.240 ;
        RECT 132.420 88.480 132.950 88.560 ;
        RECT 131.425 88.250 132.950 88.480 ;
        RECT 132.420 88.170 132.950 88.250 ;
        RECT 131.460 87.490 131.990 87.580 ;
        RECT 131.425 87.260 132.925 87.490 ;
        RECT 131.460 87.190 131.990 87.260 ;
        RECT 132.420 86.500 132.950 86.590 ;
        RECT 131.425 86.270 132.950 86.500 ;
        RECT 132.420 86.200 132.950 86.270 ;
        RECT 131.460 85.510 131.990 85.600 ;
        RECT 131.425 85.280 132.925 85.510 ;
        RECT 131.460 85.210 131.990 85.280 ;
        RECT 132.420 84.520 132.950 84.600 ;
        RECT 131.425 84.290 132.950 84.520 ;
        RECT 132.420 84.210 132.950 84.290 ;
        RECT 131.460 83.530 131.990 83.620 ;
        RECT 131.425 83.300 132.925 83.530 ;
        RECT 131.460 83.230 131.990 83.300 ;
        RECT 132.420 82.540 132.950 82.620 ;
        RECT 131.425 82.310 132.950 82.540 ;
        RECT 132.420 82.230 132.950 82.310 ;
        RECT 133.120 80.670 133.440 100.120 ;
        RECT 133.590 82.930 135.550 100.460 ;
        RECT 141.110 98.950 141.700 100.005 ;
        RECT 138.830 98.360 141.700 98.950 ;
        RECT 133.590 82.170 135.570 82.930 ;
        RECT 123.070 80.205 133.450 80.670 ;
        RECT 121.915 79.610 133.450 80.205 ;
        RECT 121.915 79.580 126.550 79.610 ;
        RECT 121.915 79.515 126.545 79.580 ;
        RECT 112.840 78.190 113.550 78.310 ;
        RECT 106.010 76.610 110.030 78.110 ;
        RECT 121.915 77.775 122.605 79.515 ;
        RECT 106.010 75.810 113.630 76.610 ;
        RECT 106.010 73.450 110.030 75.810 ;
        RECT 128.490 75.730 129.160 77.155 ;
        RECT 128.490 75.060 131.550 75.730 ;
        RECT 115.820 74.700 116.180 74.730 ;
        RECT 114.180 74.340 116.180 74.700 ;
        RECT 114.180 73.450 114.540 74.340 ;
        RECT 115.820 74.310 116.180 74.340 ;
        RECT 106.010 68.940 115.100 73.450 ;
        RECT 116.370 73.260 116.780 73.340 ;
        RECT 106.010 59.590 110.030 68.940 ;
        RECT 115.380 68.080 115.620 73.070 ;
        RECT 115.770 73.030 116.780 73.260 ;
        RECT 116.370 72.960 116.780 73.030 ;
        RECT 115.780 71.970 116.190 72.040 ;
        RECT 115.770 71.740 116.770 71.970 ;
        RECT 115.780 71.660 116.190 71.740 ;
        RECT 116.370 70.680 116.780 70.750 ;
        RECT 115.770 70.450 116.780 70.680 ;
        RECT 116.370 70.370 116.780 70.450 ;
        RECT 115.770 69.390 116.180 69.470 ;
        RECT 115.770 69.160 116.770 69.390 ;
        RECT 115.770 69.090 116.180 69.160 ;
        RECT 116.920 68.080 117.160 73.070 ;
        RECT 128.490 69.240 128.760 75.060 ;
        RECT 130.450 73.770 131.110 73.860 ;
        RECT 128.955 73.540 131.110 73.770 ;
        RECT 130.450 73.460 131.110 73.540 ;
        RECT 128.960 73.130 129.620 73.220 ;
        RECT 128.955 72.900 131.095 73.130 ;
        RECT 128.960 72.820 129.620 72.900 ;
        RECT 130.450 72.490 131.110 72.580 ;
        RECT 128.955 72.260 131.110 72.490 ;
        RECT 130.450 72.180 131.110 72.260 ;
        RECT 128.960 71.850 129.620 71.930 ;
        RECT 128.955 71.620 131.095 71.850 ;
        RECT 128.960 71.530 129.620 71.620 ;
        RECT 130.450 71.210 131.110 71.300 ;
        RECT 128.955 70.980 131.110 71.210 ;
        RECT 130.450 70.900 131.110 70.980 ;
        RECT 128.950 70.570 129.610 70.660 ;
        RECT 128.950 70.340 131.095 70.570 ;
        RECT 128.950 70.260 129.610 70.340 ;
        RECT 130.450 69.930 131.110 70.020 ;
        RECT 128.955 69.700 131.110 69.930 ;
        RECT 130.450 69.620 131.110 69.700 ;
        RECT 128.960 69.290 129.620 69.380 ;
        RECT 128.955 69.060 131.095 69.290 ;
        RECT 131.280 69.240 131.550 75.060 ;
        RECT 134.410 73.980 135.570 82.170 ;
        RECT 131.810 72.820 135.570 73.980 ;
        RECT 128.960 68.980 129.620 69.060 ;
        RECT 131.810 68.820 133.260 72.820 ;
        RECT 115.380 67.990 117.160 68.080 ;
        RECT 119.305 67.990 120.035 68.020 ;
        RECT 115.380 67.260 120.035 67.990 ;
        RECT 138.830 67.370 139.060 98.360 ;
        RECT 140.670 96.990 141.270 97.070 ;
        RECT 139.265 96.760 141.270 96.990 ;
        RECT 140.670 96.680 141.270 96.760 ;
        RECT 139.270 93.700 139.870 93.780 ;
        RECT 139.265 93.470 141.265 93.700 ;
        RECT 139.270 93.390 139.870 93.470 ;
        RECT 140.670 90.410 141.270 90.490 ;
        RECT 139.265 90.180 141.270 90.410 ;
        RECT 140.670 90.100 141.270 90.180 ;
        RECT 139.270 87.120 139.870 87.210 ;
        RECT 139.265 86.890 141.265 87.120 ;
        RECT 139.270 86.820 139.870 86.890 ;
        RECT 140.670 83.830 141.270 83.920 ;
        RECT 139.265 83.600 141.270 83.830 ;
        RECT 140.670 83.530 141.270 83.600 ;
        RECT 139.270 80.540 139.870 80.620 ;
        RECT 139.265 80.310 141.265 80.540 ;
        RECT 139.270 80.230 139.870 80.310 ;
        RECT 140.670 77.250 141.270 77.330 ;
        RECT 139.265 77.020 141.270 77.250 ;
        RECT 140.670 76.940 141.270 77.020 ;
        RECT 139.270 73.960 139.870 74.040 ;
        RECT 139.265 73.730 141.265 73.960 ;
        RECT 139.270 73.650 139.870 73.730 ;
        RECT 140.670 70.670 141.270 70.760 ;
        RECT 139.265 70.440 141.270 70.670 ;
        RECT 140.670 70.370 141.270 70.440 ;
        RECT 139.270 67.380 139.870 67.460 ;
        RECT 115.380 67.220 117.160 67.260 ;
        RECT 119.305 67.230 120.035 67.260 ;
        RECT 139.265 67.150 141.265 67.380 ;
        RECT 141.470 67.370 141.700 98.360 ;
        RECT 144.080 97.210 148.100 102.260 ;
        RECT 139.270 67.070 139.870 67.150 ;
        RECT 141.980 66.920 148.100 97.210 ;
        RECT 115.910 64.835 125.610 64.960 ;
        RECT 111.620 63.510 125.610 64.835 ;
        RECT 144.080 64.180 148.100 66.920 ;
        RECT 115.910 63.420 125.610 63.510 ;
        RECT 140.600 63.480 148.100 64.180 ;
        RECT 113.455 59.590 114.185 61.815 ;
        RECT 144.080 61.715 148.100 63.480 ;
        RECT 141.505 61.025 148.100 61.715 ;
        RECT 115.410 60.390 121.675 60.900 ;
        RECT 106.010 54.890 115.120 59.590 ;
        RECT 115.410 55.410 115.650 60.390 ;
        RECT 115.800 59.290 116.170 59.370 ;
        RECT 115.800 59.060 116.800 59.290 ;
        RECT 115.800 58.990 116.170 59.060 ;
        RECT 116.430 58.000 116.800 58.080 ;
        RECT 115.800 57.770 116.800 58.000 ;
        RECT 116.430 57.700 116.800 57.770 ;
        RECT 115.790 56.710 116.160 56.790 ;
        RECT 115.790 56.480 116.800 56.710 ;
        RECT 115.790 56.410 116.160 56.480 ;
        RECT 116.430 55.420 116.800 55.500 ;
        RECT 115.800 55.190 116.800 55.420 ;
        RECT 116.940 55.410 117.210 60.390 ;
        RECT 116.430 55.120 116.800 55.190 ;
        RECT 106.010 51.605 110.030 54.890 ;
        RECT 128.200 53.330 129.370 61.000 ;
        RECT 130.640 60.740 131.040 60.830 ;
        RECT 130.040 60.510 131.040 60.740 ;
        RECT 106.010 51.350 126.285 51.605 ;
        RECT 128.200 51.350 129.100 53.330 ;
        RECT 129.640 52.660 129.890 60.500 ;
        RECT 130.640 60.430 131.040 60.510 ;
        RECT 130.030 58.450 130.430 58.540 ;
        RECT 130.030 58.220 131.040 58.450 ;
        RECT 130.030 58.140 130.430 58.220 ;
        RECT 130.650 56.160 131.050 56.250 ;
        RECT 130.040 55.930 131.050 56.160 ;
        RECT 130.650 55.850 131.050 55.930 ;
        RECT 130.030 53.870 130.430 53.960 ;
        RECT 130.030 53.640 131.040 53.870 ;
        RECT 130.030 53.560 130.430 53.640 ;
        RECT 131.190 52.660 131.440 60.500 ;
        RECT 144.080 60.160 148.100 61.025 ;
        RECT 140.080 59.910 140.590 59.990 ;
        RECT 138.915 59.680 140.590 59.910 ;
        RECT 136.375 57.435 137.425 58.425 ;
        RECT 136.405 53.655 137.395 57.435 ;
        RECT 138.460 56.480 138.740 59.680 ;
        RECT 140.080 59.600 140.590 59.680 ;
        RECT 138.930 59.270 139.440 59.350 ;
        RECT 138.915 59.040 140.585 59.270 ;
        RECT 138.930 58.960 139.440 59.040 ;
        RECT 140.080 58.630 140.590 58.710 ;
        RECT 138.915 58.400 140.590 58.630 ;
        RECT 140.080 58.320 140.590 58.400 ;
        RECT 138.930 57.990 139.440 58.070 ;
        RECT 138.915 57.760 140.585 57.990 ;
        RECT 138.930 57.680 139.440 57.760 ;
        RECT 140.770 56.480 141.050 59.680 ;
        RECT 141.280 57.480 148.100 60.160 ;
        RECT 138.460 56.200 141.050 56.480 ;
        RECT 138.510 54.820 138.790 56.200 ;
        RECT 136.405 52.665 141.165 53.655 ;
        RECT 129.640 52.070 131.440 52.660 ;
        RECT 106.010 50.450 129.100 51.350 ;
        RECT 130.640 51.970 131.440 52.070 ;
        RECT 138.260 52.610 141.160 52.665 ;
        RECT 130.640 50.950 134.970 51.970 ;
        RECT 106.010 50.195 126.285 50.450 ;
        RECT 106.010 27.470 110.030 50.195 ;
        RECT 127.050 48.140 127.790 48.820 ;
        RECT 117.280 46.140 118.490 46.150 ;
        RECT 119.520 46.140 120.205 48.070 ;
        RECT 121.380 47.300 126.745 47.310 ;
        RECT 127.080 47.300 127.760 48.140 ;
        RECT 121.120 46.880 129.410 47.300 ;
        RECT 117.280 44.910 120.930 46.140 ;
        RECT 121.120 45.310 121.410 46.880 ;
        RECT 121.570 45.870 121.980 45.960 ;
        RECT 121.570 45.640 122.570 45.870 ;
        RECT 121.570 45.590 121.980 45.640 ;
        RECT 122.160 45.430 122.570 45.490 ;
        RECT 121.570 45.200 122.570 45.430 ;
        RECT 122.720 45.310 123.010 46.880 ;
        RECT 126.460 45.260 126.750 46.880 ;
        RECT 128.330 45.920 128.950 46.000 ;
        RECT 126.945 45.690 128.950 45.920 ;
        RECT 128.330 45.620 128.950 45.690 ;
        RECT 126.960 45.280 127.580 45.360 ;
        RECT 122.160 45.120 122.570 45.200 ;
        RECT 126.945 45.050 128.945 45.280 ;
        RECT 129.120 45.260 129.410 46.880 ;
        RECT 130.305 46.200 131.200 48.185 ;
        RECT 126.960 44.980 127.580 45.050 ;
        RECT 117.280 41.460 120.060 44.910 ;
        RECT 129.630 44.790 132.730 46.200 ;
        RECT 124.480 43.260 125.165 44.435 ;
        RECT 121.380 43.250 129.420 43.260 ;
        RECT 121.150 42.820 129.420 43.250 ;
        RECT 121.150 42.800 126.750 42.820 ;
        RECT 117.280 39.750 120.910 41.460 ;
        RECT 121.150 40.640 121.430 42.800 ;
        RECT 122.600 41.190 123.030 41.270 ;
        RECT 121.570 40.960 123.070 41.190 ;
        RECT 122.600 40.870 123.030 40.960 ;
        RECT 121.620 40.710 122.050 40.790 ;
        RECT 121.570 40.480 123.070 40.710 ;
        RECT 121.620 40.390 122.050 40.480 ;
        RECT 122.600 40.230 123.030 40.320 ;
        RECT 121.570 40.000 123.070 40.230 ;
        RECT 123.210 40.160 123.500 42.800 ;
        RECT 122.600 39.920 123.030 40.000 ;
        RECT 126.460 39.870 126.740 42.800 ;
        RECT 128.380 41.780 128.940 41.870 ;
        RECT 126.945 41.550 128.945 41.780 ;
        RECT 128.380 41.470 128.940 41.550 ;
        RECT 126.960 41.140 127.520 41.220 ;
        RECT 126.945 40.910 128.945 41.140 ;
        RECT 126.960 40.820 127.520 40.910 ;
        RECT 128.380 40.500 128.940 40.590 ;
        RECT 126.945 40.270 128.945 40.500 ;
        RECT 128.380 40.190 128.940 40.270 ;
        RECT 126.960 39.860 127.520 39.940 ;
        RECT 129.130 39.870 129.410 42.820 ;
        RECT 130.810 42.050 132.730 44.790 ;
        RECT 117.280 34.620 118.490 39.750 ;
        RECT 126.945 39.630 128.945 39.860 ;
        RECT 126.960 39.540 127.520 39.630 ;
        RECT 129.620 39.360 132.730 42.050 ;
        RECT 119.510 37.560 121.900 38.240 ;
        RECT 124.405 37.560 125.280 39.060 ;
        RECT 119.510 37.540 126.865 37.560 ;
        RECT 119.510 36.870 130.400 37.540 ;
        RECT 119.510 36.850 126.865 36.870 ;
        RECT 119.510 36.695 121.900 36.850 ;
        RECT 117.280 32.430 119.470 34.620 ;
        RECT 119.710 32.860 119.980 36.695 ;
        RECT 120.190 34.360 120.700 34.460 ;
        RECT 120.130 34.130 123.130 34.360 ;
        RECT 120.190 34.030 120.700 34.130 ;
        RECT 122.570 33.880 123.080 33.980 ;
        RECT 120.130 33.650 123.130 33.880 ;
        RECT 122.570 33.550 123.080 33.650 ;
        RECT 120.200 33.400 120.710 33.500 ;
        RECT 120.130 33.170 123.130 33.400 ;
        RECT 123.280 33.340 123.550 36.850 ;
        RECT 120.200 33.070 120.710 33.170 ;
        RECT 122.570 32.920 123.080 33.020 ;
        RECT 120.130 32.690 123.130 32.920 ;
        RECT 122.570 32.590 123.080 32.690 ;
        RECT 117.280 27.470 118.940 32.430 ;
        RECT 126.460 31.700 126.740 36.850 ;
        RECT 129.340 35.560 129.940 35.640 ;
        RECT 126.945 35.330 129.945 35.560 ;
        RECT 129.340 35.240 129.940 35.330 ;
        RECT 126.980 34.920 127.580 35.000 ;
        RECT 126.945 34.690 129.945 34.920 ;
        RECT 126.980 34.600 127.580 34.690 ;
        RECT 129.340 34.280 129.940 34.370 ;
        RECT 126.945 34.050 129.945 34.280 ;
        RECT 129.340 33.970 129.940 34.050 ;
        RECT 126.980 33.640 127.580 33.730 ;
        RECT 126.945 33.410 129.945 33.640 ;
        RECT 126.980 33.330 127.580 33.410 ;
        RECT 129.340 33.000 129.940 33.080 ;
        RECT 126.945 32.770 129.945 33.000 ;
        RECT 129.340 32.680 129.940 32.770 ;
        RECT 126.980 32.360 127.580 32.450 ;
        RECT 126.945 32.130 129.945 32.360 ;
        RECT 126.980 32.050 127.580 32.130 ;
        RECT 129.340 31.720 129.940 31.810 ;
        RECT 126.945 31.490 129.945 31.720 ;
        RECT 130.120 31.700 130.400 36.870 ;
        RECT 131.580 35.760 132.730 39.360 ;
        RECT 129.340 31.410 129.940 31.490 ;
        RECT 130.650 31.240 132.730 35.760 ;
        RECT 133.950 34.395 134.970 50.950 ;
        RECT 106.010 25.810 118.940 27.470 ;
        RECT 123.960 27.125 125.040 29.540 ;
        RECT 130.920 27.295 132.730 31.240 ;
        RECT 133.845 29.495 135.015 34.395 ;
        RECT 138.260 31.600 138.520 52.610 ;
        RECT 138.730 51.350 139.300 51.450 ;
        RECT 138.715 51.120 140.715 51.350 ;
        RECT 138.730 51.030 139.300 51.120 ;
        RECT 140.150 48.060 140.720 48.160 ;
        RECT 138.715 47.830 140.720 48.060 ;
        RECT 140.150 47.740 140.720 47.830 ;
        RECT 138.730 44.770 139.300 44.880 ;
        RECT 138.715 44.540 140.715 44.770 ;
        RECT 138.730 44.460 139.300 44.540 ;
        RECT 140.160 41.480 140.730 41.580 ;
        RECT 138.715 41.250 140.730 41.480 ;
        RECT 140.160 41.160 140.730 41.250 ;
        RECT 138.730 38.190 139.300 38.290 ;
        RECT 138.715 37.960 140.715 38.190 ;
        RECT 138.730 37.870 139.300 37.960 ;
        RECT 140.160 34.900 140.730 35.000 ;
        RECT 138.715 34.670 140.730 34.900 ;
        RECT 140.160 34.580 140.730 34.670 ;
        RECT 138.730 31.610 139.300 31.700 ;
        RECT 138.715 31.380 140.715 31.610 ;
        RECT 140.900 31.600 141.160 52.610 ;
        RECT 144.080 51.610 148.100 57.480 ;
        RECT 138.730 31.280 139.300 31.380 ;
        RECT 141.440 31.080 148.100 51.610 ;
        RECT 144.080 29.575 148.100 31.080 ;
        RECT 140.035 28.760 148.100 29.575 ;
        RECT 144.080 27.295 148.100 28.760 ;
        RECT 106.010 25.010 110.030 25.810 ;
        RECT 123.875 19.435 125.045 27.125 ;
        RECT 130.920 25.485 148.100 27.295 ;
        RECT 144.080 25.010 148.100 25.485 ;
      LAYER via ;
        RECT 145.140 141.540 146.640 143.040 ;
        RECT 137.000 129.090 137.600 129.690 ;
        RECT 118.970 113.940 119.530 114.500 ;
        RECT 124.310 118.900 124.800 119.190 ;
        RECT 121.870 118.440 122.360 118.730 ;
        RECT 124.310 117.960 124.800 118.250 ;
        RECT 121.870 117.480 122.360 117.770 ;
        RECT 124.310 117.000 124.800 117.290 ;
        RECT 121.870 116.520 122.360 116.810 ;
        RECT 124.310 116.040 124.800 116.330 ;
        RECT 121.870 115.560 122.360 115.850 ;
        RECT 123.495 113.990 124.065 114.560 ;
        RECT 127.230 115.430 128.795 116.995 ;
        RECT 131.050 118.860 131.530 119.140 ;
        RECT 133.450 118.290 133.930 118.570 ;
        RECT 131.030 117.640 131.510 117.920 ;
        RECT 133.450 117.000 133.930 117.280 ;
        RECT 131.030 116.370 131.510 116.650 ;
        RECT 133.450 115.730 133.930 116.010 ;
        RECT 131.030 115.080 131.510 115.360 ;
        RECT 133.450 114.450 133.930 114.730 ;
        RECT 131.000 112.730 131.580 113.310 ;
        RECT 141.110 109.775 141.700 110.365 ;
        RECT 116.020 103.730 116.650 104.050 ;
        RECT 112.790 100.460 113.420 100.780 ;
        RECT 116.020 97.150 116.650 97.470 ;
        RECT 112.790 93.850 113.420 94.170 ;
        RECT 112.740 91.790 113.490 92.540 ;
        RECT 116.020 88.100 116.730 88.470 ;
        RECT 112.840 84.810 113.550 85.180 ;
        RECT 116.020 81.530 116.730 81.900 ;
        RECT 112.840 78.240 113.550 78.610 ;
        RECT 124.630 100.100 125.040 100.390 ;
        RECT 123.650 99.110 124.060 99.400 ;
        RECT 124.630 98.120 125.040 98.410 ;
        RECT 123.650 97.130 124.060 97.420 ;
        RECT 124.630 96.140 125.040 96.430 ;
        RECT 123.650 95.150 124.060 95.440 ;
        RECT 124.630 94.160 125.040 94.450 ;
        RECT 123.650 93.180 124.060 93.470 ;
        RECT 124.630 92.180 125.040 92.470 ;
        RECT 123.650 91.200 124.060 91.490 ;
        RECT 124.630 90.200 125.040 90.490 ;
        RECT 123.650 89.210 124.060 89.500 ;
        RECT 124.630 88.220 125.040 88.510 ;
        RECT 123.650 87.240 124.060 87.530 ;
        RECT 124.630 86.240 125.040 86.530 ;
        RECT 123.650 85.250 124.060 85.540 ;
        RECT 124.630 84.260 125.040 84.550 ;
        RECT 123.650 83.270 124.060 83.560 ;
        RECT 124.630 82.280 125.040 82.570 ;
        RECT 132.420 100.100 132.950 100.390 ;
        RECT 131.460 99.110 131.990 99.400 ;
        RECT 132.420 98.120 132.950 98.410 ;
        RECT 131.460 97.140 131.990 97.430 ;
        RECT 132.420 96.140 132.950 96.430 ;
        RECT 131.460 95.160 131.990 95.450 ;
        RECT 132.420 94.170 132.950 94.460 ;
        RECT 131.460 93.170 131.990 93.460 ;
        RECT 132.420 92.190 132.950 92.480 ;
        RECT 131.460 91.190 131.990 91.480 ;
        RECT 132.420 90.200 132.950 90.490 ;
        RECT 131.460 89.220 131.990 89.510 ;
        RECT 132.420 88.220 132.950 88.510 ;
        RECT 131.460 87.240 131.990 87.530 ;
        RECT 132.420 86.250 132.950 86.540 ;
        RECT 131.460 85.260 131.990 85.550 ;
        RECT 132.420 84.260 132.950 84.550 ;
        RECT 131.460 83.280 131.990 83.570 ;
        RECT 132.420 82.280 132.950 82.570 ;
        RECT 141.110 99.385 141.700 99.975 ;
        RECT 121.915 77.805 122.605 78.495 ;
        RECT 112.800 75.810 113.600 76.610 ;
        RECT 128.490 76.455 129.160 77.125 ;
        RECT 115.820 74.340 116.180 74.700 ;
        RECT 116.370 73.010 116.780 73.290 ;
        RECT 115.780 71.710 116.190 71.990 ;
        RECT 116.370 70.420 116.780 70.700 ;
        RECT 115.770 69.140 116.180 69.420 ;
        RECT 130.450 73.510 131.110 73.810 ;
        RECT 128.960 72.870 129.620 73.170 ;
        RECT 130.450 72.230 131.110 72.530 ;
        RECT 128.960 71.580 129.620 71.880 ;
        RECT 130.450 70.950 131.110 71.250 ;
        RECT 128.950 70.310 129.610 70.610 ;
        RECT 130.450 69.670 131.110 69.970 ;
        RECT 128.960 69.030 129.620 69.330 ;
        RECT 116.430 67.535 116.820 67.925 ;
        RECT 119.305 67.260 120.035 67.990 ;
        RECT 140.670 96.730 141.270 97.020 ;
        RECT 139.270 93.440 139.870 93.730 ;
        RECT 140.670 90.150 141.270 90.440 ;
        RECT 139.270 86.870 139.870 87.160 ;
        RECT 140.670 83.580 141.270 83.870 ;
        RECT 139.270 80.280 139.870 80.570 ;
        RECT 140.670 76.990 141.270 77.280 ;
        RECT 139.270 73.700 139.870 73.990 ;
        RECT 140.670 70.420 141.270 70.710 ;
        RECT 139.270 67.120 139.870 67.410 ;
        RECT 111.980 63.870 112.580 64.470 ;
        RECT 124.040 63.420 125.580 64.960 ;
        RECT 140.630 63.480 141.330 64.180 ;
        RECT 113.455 61.055 114.185 61.785 ;
        RECT 141.560 61.080 142.140 61.660 ;
        RECT 121.135 60.390 121.645 60.900 ;
        RECT 115.800 59.040 116.170 59.320 ;
        RECT 116.430 57.750 116.800 58.030 ;
        RECT 115.790 56.460 116.160 56.740 ;
        RECT 116.430 55.170 116.800 55.450 ;
        RECT 130.640 60.480 131.040 60.780 ;
        RECT 130.030 58.190 130.430 58.490 ;
        RECT 130.650 55.900 131.050 56.200 ;
        RECT 130.030 53.610 130.430 53.910 ;
        RECT 136.405 57.435 137.395 58.425 ;
        RECT 140.080 59.650 140.590 59.940 ;
        RECT 138.930 59.010 139.440 59.300 ;
        RECT 140.080 58.370 140.590 58.660 ;
        RECT 138.930 57.730 139.440 58.020 ;
        RECT 138.510 54.850 138.790 55.130 ;
        RECT 127.080 48.140 127.760 48.820 ;
        RECT 119.605 47.475 120.115 47.985 ;
        RECT 130.385 47.375 131.115 48.105 ;
        RECT 122.160 45.170 122.570 45.440 ;
        RECT 128.330 45.670 128.950 45.950 ;
        RECT 126.960 45.030 127.580 45.310 ;
        RECT 124.555 43.830 125.085 44.360 ;
        RECT 118.910 42.000 119.430 42.520 ;
        RECT 131.215 42.945 131.865 43.595 ;
        RECT 122.600 40.920 123.030 41.220 ;
        RECT 121.620 40.440 122.050 40.740 ;
        RECT 122.600 39.970 123.030 40.270 ;
        RECT 128.380 41.520 128.940 41.820 ;
        RECT 126.960 40.870 127.520 41.170 ;
        RECT 128.380 40.240 128.940 40.540 ;
        RECT 126.960 39.590 127.520 39.890 ;
        RECT 124.515 38.300 125.165 38.950 ;
        RECT 119.715 36.905 120.845 38.035 ;
        RECT 120.190 34.080 120.700 34.410 ;
        RECT 122.570 33.600 123.080 33.930 ;
        RECT 120.200 33.120 120.710 33.450 ;
        RECT 122.570 32.640 123.080 32.970 ;
        RECT 129.340 35.290 129.940 35.590 ;
        RECT 126.980 34.650 127.580 34.950 ;
        RECT 129.340 34.020 129.940 34.320 ;
        RECT 126.980 33.380 127.580 33.680 ;
        RECT 129.340 32.730 129.940 33.030 ;
        RECT 126.980 32.100 127.580 32.400 ;
        RECT 129.340 31.460 129.940 31.760 ;
        RECT 117.925 30.600 118.555 31.230 ;
        RECT 131.335 29.620 132.105 30.390 ;
        RECT 124.185 28.685 124.815 29.315 ;
        RECT 138.730 51.080 139.300 51.400 ;
        RECT 140.150 47.790 140.720 48.110 ;
        RECT 138.730 44.510 139.300 44.830 ;
        RECT 140.160 41.210 140.730 41.530 ;
        RECT 138.730 37.920 139.300 38.240 ;
        RECT 140.160 34.630 140.730 34.950 ;
        RECT 138.730 31.330 139.300 31.650 ;
        RECT 134.130 29.780 134.730 30.380 ;
        RECT 140.120 28.850 140.760 29.490 ;
        RECT 124.160 19.720 124.760 20.320 ;
      LAYER met2 ;
        RECT 96.485 143.040 97.935 143.060 ;
        RECT 96.460 141.540 146.670 143.040 ;
        RECT 96.485 141.520 97.935 141.540 ;
        RECT 76.935 134.210 78.385 134.230 ;
        RECT 76.910 132.710 88.430 134.210 ;
        RECT 76.935 132.690 78.385 132.710 ;
        RECT 136.970 129.090 157.160 129.690 ;
        RECT 124.260 118.900 124.850 119.190 ;
        RECT 121.820 118.440 122.410 118.730 ;
        RECT 121.850 117.770 122.410 118.440 ;
        RECT 124.280 118.250 124.850 118.900 ;
        RECT 124.260 117.960 124.850 118.250 ;
        RECT 121.820 117.480 122.410 117.770 ;
        RECT 121.850 116.810 122.410 117.480 ;
        RECT 124.280 117.290 124.850 117.960 ;
        RECT 131.000 117.920 131.580 119.150 ;
        RECT 133.420 118.570 133.960 118.630 ;
        RECT 133.400 118.290 133.980 118.570 ;
        RECT 130.980 117.640 131.580 117.920 ;
        RECT 124.260 117.000 124.850 117.290 ;
        RECT 121.820 116.520 122.410 116.810 ;
        RECT 121.850 115.850 122.410 116.520 ;
        RECT 124.280 116.330 124.850 117.000 ;
        RECT 124.260 116.040 124.850 116.330 ;
        RECT 121.820 115.560 122.410 115.850 ;
        RECT 118.970 114.500 119.530 114.530 ;
        RECT 121.850 114.500 122.410 115.560 ;
        RECT 124.280 114.560 124.850 116.040 ;
        RECT 127.200 115.430 128.825 116.995 ;
        RECT 131.000 116.650 131.580 117.640 ;
        RECT 133.420 117.280 133.960 118.290 ;
        RECT 133.400 117.000 133.980 117.280 ;
        RECT 130.980 116.370 131.580 116.650 ;
        RECT 118.970 113.940 122.410 114.500 ;
        RECT 123.465 113.990 124.850 114.560 ;
        RECT 118.970 113.910 119.530 113.940 ;
        RECT 127.230 107.785 128.795 115.430 ;
        RECT 131.000 115.360 131.580 116.370 ;
        RECT 133.420 116.010 133.960 117.000 ;
        RECT 133.400 115.730 133.980 116.010 ;
        RECT 130.980 115.080 131.580 115.360 ;
        RECT 131.000 112.700 131.580 115.080 ;
        RECT 133.420 114.730 133.960 115.730 ;
        RECT 133.400 114.450 133.980 114.730 ;
        RECT 133.420 113.270 133.960 114.450 ;
        RECT 133.420 112.730 136.490 113.270 ;
        RECT 115.970 105.580 125.185 106.290 ;
        RECT 127.230 106.220 133.440 107.785 ;
        RECT 115.970 104.050 116.680 105.580 ;
        RECT 115.970 103.730 116.700 104.050 ;
        RECT 112.740 91.760 113.490 100.850 ;
        RECT 115.970 97.470 116.680 103.730 ;
        RECT 124.475 103.205 125.185 105.580 ;
        RECT 131.875 104.070 133.440 106.220 ;
        RECT 131.420 103.205 132.010 103.230 ;
        RECT 124.475 102.495 132.010 103.205 ;
        RECT 124.590 100.390 125.100 100.440 ;
        RECT 124.580 100.100 125.100 100.390 ;
        RECT 115.970 97.150 116.700 97.470 ;
        RECT 115.970 96.750 116.680 97.150 ;
        RECT 115.950 88.470 116.750 88.580 ;
        RECT 115.950 88.100 116.780 88.470 ;
        RECT 112.800 85.180 113.600 85.290 ;
        RECT 112.790 84.810 113.600 85.180 ;
        RECT 112.800 78.610 113.600 84.810 ;
        RECT 112.790 78.240 113.600 78.610 ;
        RECT 112.800 75.780 113.600 78.240 ;
        RECT 115.950 81.900 116.750 88.100 ;
        RECT 115.950 81.530 116.780 81.900 ;
        RECT 115.950 76.800 116.750 81.530 ;
        RECT 123.540 78.660 124.200 99.600 ;
        RECT 124.590 98.410 125.100 100.100 ;
        RECT 124.580 98.120 125.100 98.410 ;
        RECT 124.590 96.430 125.100 98.120 ;
        RECT 124.580 96.140 125.100 96.430 ;
        RECT 124.590 94.450 125.100 96.140 ;
        RECT 124.580 94.160 125.100 94.450 ;
        RECT 124.590 92.470 125.100 94.160 ;
        RECT 124.580 92.180 125.100 92.470 ;
        RECT 124.590 90.490 125.100 92.180 ;
        RECT 124.580 90.200 125.100 90.490 ;
        RECT 124.590 88.510 125.100 90.200 ;
        RECT 124.580 88.220 125.100 88.510 ;
        RECT 124.590 86.530 125.100 88.220 ;
        RECT 124.580 86.240 125.100 86.530 ;
        RECT 124.590 84.550 125.100 86.240 ;
        RECT 124.580 84.260 125.100 84.550 ;
        RECT 124.590 82.570 125.100 84.260 ;
        RECT 124.580 82.280 125.100 82.570 ;
        RECT 123.540 78.495 124.230 78.660 ;
        RECT 121.885 77.805 124.230 78.495 ;
        RECT 123.540 77.600 124.230 77.805 ;
        RECT 123.540 76.800 124.200 77.600 ;
        RECT 115.950 76.000 124.270 76.800 ;
        RECT 124.590 75.595 125.100 82.280 ;
        RECT 128.490 77.125 129.160 102.495 ;
        RECT 131.420 99.400 132.010 102.495 ;
        RECT 132.320 100.390 132.990 104.070 ;
        RECT 136.405 101.015 137.395 101.215 ;
        RECT 141.110 101.015 141.700 110.395 ;
        RECT 156.560 102.985 157.160 129.090 ;
        RECT 156.540 102.435 157.180 102.985 ;
        RECT 156.560 102.410 157.160 102.435 ;
        RECT 136.405 100.425 141.700 101.015 ;
        RECT 132.320 100.100 133.000 100.390 ;
        RECT 131.410 99.110 132.040 99.400 ;
        RECT 131.420 97.430 132.010 99.110 ;
        RECT 132.320 98.410 132.990 100.100 ;
        RECT 132.320 98.120 133.000 98.410 ;
        RECT 131.410 97.140 132.040 97.430 ;
        RECT 131.420 95.450 132.010 97.140 ;
        RECT 132.320 96.430 132.990 98.120 ;
        RECT 132.320 96.140 133.000 96.430 ;
        RECT 131.410 95.160 132.040 95.450 ;
        RECT 131.420 93.460 132.010 95.160 ;
        RECT 132.320 94.460 132.990 96.140 ;
        RECT 132.320 94.170 133.000 94.460 ;
        RECT 131.410 93.170 132.040 93.460 ;
        RECT 131.420 91.480 132.010 93.170 ;
        RECT 132.320 92.480 132.990 94.170 ;
        RECT 132.320 92.190 133.000 92.480 ;
        RECT 131.410 91.190 132.040 91.480 ;
        RECT 131.420 89.510 132.010 91.190 ;
        RECT 132.320 90.490 132.990 92.190 ;
        RECT 132.320 90.200 133.000 90.490 ;
        RECT 131.410 89.220 132.040 89.510 ;
        RECT 131.420 87.530 132.010 89.220 ;
        RECT 132.320 88.510 132.990 90.200 ;
        RECT 132.320 88.220 133.000 88.510 ;
        RECT 131.410 87.240 132.040 87.530 ;
        RECT 131.420 85.550 132.010 87.240 ;
        RECT 132.320 86.540 132.990 88.220 ;
        RECT 132.320 86.250 133.000 86.540 ;
        RECT 131.410 85.260 132.040 85.550 ;
        RECT 131.420 83.570 132.010 85.260 ;
        RECT 132.320 84.550 132.990 86.250 ;
        RECT 132.320 84.260 133.000 84.550 ;
        RECT 131.410 83.280 132.040 83.570 ;
        RECT 131.420 83.160 132.010 83.280 ;
        RECT 132.320 82.570 132.990 84.260 ;
        RECT 132.320 82.280 133.000 82.570 ;
        RECT 132.320 82.245 132.990 82.280 ;
        RECT 128.460 76.455 129.190 77.125 ;
        RECT 124.590 75.085 134.885 75.595 ;
        RECT 115.790 74.340 116.210 74.700 ;
        RECT 115.820 71.990 116.180 74.340 ;
        RECT 116.320 73.010 116.830 73.290 ;
        RECT 128.970 73.170 129.700 73.220 ;
        RECT 115.730 71.710 116.240 71.990 ;
        RECT 115.820 69.420 116.180 71.710 ;
        RECT 116.430 70.700 116.820 73.010 ;
        RECT 128.910 72.870 129.700 73.170 ;
        RECT 128.970 71.880 129.700 72.870 ;
        RECT 128.910 71.580 129.700 71.880 ;
        RECT 116.320 70.420 116.830 70.700 ;
        RECT 128.970 70.610 129.700 71.580 ;
        RECT 115.720 69.140 116.230 69.420 ;
        RECT 115.820 69.130 116.180 69.140 ;
        RECT 116.430 67.505 116.820 70.420 ;
        RECT 128.900 70.310 129.700 70.610 ;
        RECT 128.970 69.330 129.700 70.310 ;
        RECT 130.390 69.520 131.160 75.085 ;
        RECT 128.910 69.030 129.700 69.330 ;
        RECT 128.970 67.990 129.700 69.030 ;
        RECT 119.275 67.260 129.700 67.990 ;
        RECT 90.320 63.870 112.610 64.470 ;
        RECT 90.320 37.405 90.920 63.870 ;
        RECT 113.425 61.650 114.895 61.785 ;
        RECT 113.425 61.190 116.210 61.650 ;
        RECT 113.425 61.055 114.895 61.190 ;
        RECT 115.750 59.320 116.210 61.190 ;
        RECT 120.990 60.240 121.795 67.260 ;
        RECT 134.375 66.825 134.885 75.085 ;
        RECT 136.405 68.740 137.395 100.425 ;
        RECT 141.110 99.975 141.700 100.425 ;
        RECT 141.080 99.385 141.730 99.975 ;
        RECT 140.630 97.020 141.330 97.080 ;
        RECT 140.620 96.730 141.330 97.020 ;
        RECT 139.230 93.730 139.930 93.830 ;
        RECT 139.220 93.440 139.930 93.730 ;
        RECT 139.230 87.160 139.930 93.440 ;
        RECT 140.630 90.440 141.330 96.730 ;
        RECT 140.620 90.150 141.330 90.440 ;
        RECT 139.220 86.870 139.930 87.160 ;
        RECT 139.230 80.570 139.930 86.870 ;
        RECT 140.630 83.870 141.330 90.150 ;
        RECT 140.620 83.580 141.330 83.870 ;
        RECT 139.220 80.280 139.930 80.570 ;
        RECT 139.230 73.990 139.930 80.280 ;
        RECT 140.630 77.280 141.330 83.580 ;
        RECT 140.620 76.990 141.330 77.280 ;
        RECT 139.220 73.700 139.930 73.990 ;
        RECT 139.230 67.410 139.930 73.700 ;
        RECT 140.630 70.710 141.330 76.990 ;
        RECT 140.620 70.420 141.330 70.710 ;
        RECT 139.220 67.120 139.930 67.410 ;
        RECT 134.365 66.255 134.885 66.825 ;
        RECT 134.365 65.320 134.875 66.255 ;
        RECT 139.230 65.320 139.930 67.120 ;
        RECT 124.040 64.960 125.580 64.990 ;
        RECT 124.040 64.930 130.450 64.960 ;
        RECT 134.360 64.930 139.930 65.320 ;
        RECT 124.040 63.485 139.930 64.930 ;
        RECT 124.040 63.420 130.450 63.485 ;
        RECT 134.360 63.480 139.930 63.485 ;
        RECT 140.630 63.450 141.330 70.420 ;
        RECT 124.040 63.390 125.580 63.420 ;
        RECT 115.750 59.040 116.220 59.320 ;
        RECT 115.750 56.740 116.210 59.040 ;
        RECT 129.970 58.490 130.430 63.420 ;
        RECT 130.640 61.690 139.480 62.140 ;
        RECT 130.640 60.780 131.090 61.690 ;
        RECT 130.590 60.480 131.090 60.780 ;
        RECT 129.970 58.190 130.480 58.490 ;
        RECT 116.400 58.030 116.850 58.060 ;
        RECT 116.380 57.750 116.850 58.030 ;
        RECT 115.740 56.460 116.210 56.740 ;
        RECT 115.750 56.430 116.210 56.460 ;
        RECT 116.400 55.450 116.850 57.750 ;
        RECT 116.380 55.170 116.850 55.450 ;
        RECT 116.400 53.390 116.850 55.170 ;
        RECT 129.970 53.910 130.430 58.190 ;
        RECT 130.640 56.200 131.090 60.480 ;
        RECT 136.405 59.870 137.395 59.895 ;
        RECT 130.600 55.900 131.100 56.200 ;
        RECT 133.825 55.975 134.955 59.860 ;
        RECT 136.385 58.930 137.415 59.870 ;
        RECT 138.870 59.300 139.480 61.690 ;
        RECT 140.060 61.080 142.170 61.660 ;
        RECT 140.060 59.940 140.640 61.080 ;
        RECT 140.030 59.650 140.640 59.940 ;
        RECT 138.870 59.010 139.490 59.300 ;
        RECT 136.405 57.405 137.395 58.930 ;
        RECT 138.870 58.020 139.480 59.010 ;
        RECT 140.060 58.660 140.640 59.650 ;
        RECT 140.030 58.370 140.640 58.660 ;
        RECT 140.060 58.330 140.640 58.370 ;
        RECT 138.870 57.730 139.490 58.020 ;
        RECT 138.870 57.710 139.480 57.730 ;
        RECT 130.640 55.800 131.090 55.900 ;
        RECT 134.080 55.300 134.705 55.975 ;
        RECT 134.080 54.675 138.965 55.300 ;
        RECT 129.970 53.610 130.480 53.910 ;
        RECT 129.970 53.570 130.430 53.610 ;
        RECT 116.400 52.125 127.760 53.390 ;
        RECT 116.780 52.100 127.760 52.125 ;
        RECT 127.070 50.040 127.750 52.100 ;
        RECT 127.070 49.450 132.610 50.040 ;
        RECT 127.070 49.435 135.210 49.450 ;
        RECT 127.070 49.360 137.205 49.435 ;
        RECT 127.080 48.110 127.760 49.360 ;
        RECT 131.930 48.770 137.205 49.360 ;
        RECT 134.665 48.745 137.205 48.770 ;
        RECT 119.575 47.475 122.030 47.985 ;
        RECT 121.520 45.640 122.030 47.475 ;
        RECT 128.280 47.375 131.145 48.105 ;
        RECT 128.280 45.670 129.010 47.375 ;
        RECT 122.110 44.360 122.640 45.440 ;
        RECT 126.900 44.360 127.630 45.320 ;
        RECT 122.110 43.830 127.630 44.360 ;
        RECT 128.340 42.945 131.895 43.595 ;
        RECT 118.880 42.000 122.090 42.520 ;
        RECT 121.570 40.740 122.090 42.000 ;
        RECT 128.340 41.820 128.990 42.945 ;
        RECT 128.330 41.520 128.990 41.820 ;
        RECT 122.580 41.220 123.080 41.240 ;
        RECT 122.550 40.920 123.080 41.220 ;
        RECT 121.570 40.440 122.100 40.740 ;
        RECT 121.570 40.410 122.090 40.440 ;
        RECT 122.580 40.270 123.080 40.920 ;
        RECT 122.550 39.970 123.080 40.270 ;
        RECT 122.580 38.950 123.080 39.970 ;
        RECT 126.910 41.170 127.560 41.210 ;
        RECT 126.910 40.870 127.570 41.170 ;
        RECT 126.910 39.890 127.560 40.870 ;
        RECT 128.340 40.540 128.990 41.520 ;
        RECT 128.330 40.240 128.990 40.540 ;
        RECT 128.340 40.220 128.990 40.240 ;
        RECT 126.910 39.590 127.570 39.890 ;
        RECT 124.515 38.950 125.165 38.980 ;
        RECT 126.910 38.950 127.560 39.590 ;
        RECT 122.575 38.300 127.560 38.950 ;
        RECT 122.580 38.280 123.080 38.300 ;
        RECT 124.515 38.270 125.165 38.300 ;
        RECT 114.055 38.010 120.875 38.035 ;
        RECT 90.300 36.855 90.940 37.405 ;
        RECT 114.035 36.930 120.875 38.010 ;
        RECT 114.055 36.905 120.875 36.930 ;
        RECT 90.320 36.830 90.920 36.855 ;
        RECT 120.130 31.230 120.760 34.460 ;
        RECT 117.895 30.600 120.760 31.230 ;
        RECT 122.500 30.240 123.130 33.940 ;
        RECT 126.930 30.240 127.640 34.960 ;
        RECT 122.500 29.610 127.640 30.240 ;
        RECT 129.230 30.390 130.000 35.650 ;
        RECT 129.230 29.620 132.135 30.390 ;
        RECT 124.185 28.655 124.815 29.610 ;
        RECT 134.130 28.930 134.730 30.410 ;
        RECT 136.515 30.220 137.205 48.745 ;
        RECT 138.660 30.220 139.350 51.460 ;
        RECT 140.120 48.110 140.760 48.200 ;
        RECT 140.100 47.790 140.770 48.110 ;
        RECT 140.120 41.530 140.760 47.790 ;
        RECT 140.110 41.210 140.780 41.530 ;
        RECT 140.120 34.950 140.760 41.210 ;
        RECT 140.110 34.630 140.780 34.950 ;
        RECT 136.515 29.530 139.350 30.220 ;
        RECT 140.120 29.490 140.760 34.630 ;
        RECT 134.130 28.330 135.080 28.930 ;
        RECT 140.090 28.850 140.790 29.490 ;
        RECT 124.160 12.905 124.760 20.350 ;
        RECT 134.480 15.955 135.080 28.330 ;
        RECT 134.460 15.405 135.100 15.955 ;
        RECT 134.480 15.380 135.080 15.405 ;
        RECT 124.140 12.355 124.780 12.905 ;
        RECT 124.160 12.330 124.760 12.355 ;
      LAYER via2 ;
        RECT 96.485 141.565 97.935 143.015 ;
        RECT 76.935 132.735 78.385 134.185 ;
        RECT 156.585 102.435 157.135 102.985 ;
        RECT 136.405 68.785 137.395 69.775 ;
        RECT 133.825 58.685 134.955 59.815 ;
        RECT 136.430 58.930 137.370 59.870 ;
        RECT 90.345 36.855 90.895 37.405 ;
        RECT 114.080 36.930 115.160 38.010 ;
        RECT 134.505 15.405 135.055 15.955 ;
        RECT 124.185 12.355 124.735 12.905 ;
      LAYER met3 ;
        RECT 29.685 143.040 31.175 143.065 ;
        RECT 29.680 141.540 97.960 143.040 ;
        RECT 29.685 141.515 31.175 141.540 ;
        RECT 69.815 134.210 71.305 134.235 ;
        RECT 69.810 132.710 78.410 134.210 ;
        RECT 69.815 132.685 71.305 132.710 ;
        RECT 136.380 68.760 137.420 69.800 ;
        RECT 126.305 62.565 134.955 63.695 ;
        RECT 126.305 56.955 127.435 62.565 ;
        RECT 133.825 59.840 134.955 62.565 ;
        RECT 133.800 58.660 134.980 59.840 ;
        RECT 136.405 58.905 137.395 68.760 ;
        RECT 120.335 55.825 127.435 56.955 ;
        RECT 120.335 51.055 121.465 55.825 ;
        RECT 114.055 49.925 121.465 51.055 ;
        RECT 90.320 22.915 90.920 37.430 ;
        RECT 114.055 36.905 115.185 49.925 ;
        RECT 156.560 47.445 157.160 103.010 ;
        RECT 156.535 46.855 157.185 47.445 ;
        RECT 156.560 46.850 157.160 46.855 ;
        RECT 90.295 22.325 90.945 22.915 ;
        RECT 90.320 22.320 90.920 22.325 ;
        RECT 117.785 11.050 118.375 11.075 ;
        RECT 124.160 11.050 124.760 12.930 ;
        RECT 134.480 11.265 135.080 15.980 ;
        RECT 117.780 10.450 124.760 11.050 ;
        RECT 134.455 10.675 135.105 11.265 ;
        RECT 134.480 10.670 135.080 10.675 ;
        RECT 117.785 10.425 118.375 10.450 ;
      LAYER via3 ;
        RECT 29.685 141.545 31.175 143.035 ;
        RECT 69.815 132.715 71.305 134.205 ;
        RECT 156.565 46.855 157.155 47.445 ;
        RECT 90.325 22.325 90.915 22.915 ;
        RECT 117.785 10.455 118.375 11.045 ;
        RECT 134.485 10.675 135.075 11.265 ;
      LAYER met4 ;
        RECT 3.990 224.190 4.290 224.760 ;
        RECT 7.670 224.190 7.970 224.760 ;
        RECT 11.350 224.190 11.650 224.760 ;
        RECT 15.030 224.190 15.330 224.760 ;
        RECT 18.710 224.190 19.010 224.760 ;
        RECT 22.390 224.190 22.690 224.760 ;
        RECT 26.070 224.190 26.370 224.760 ;
        RECT 29.750 224.190 30.050 224.760 ;
        RECT 33.430 224.190 33.730 224.760 ;
        RECT 37.110 224.190 37.410 224.760 ;
        RECT 40.790 224.190 41.090 224.760 ;
        RECT 44.470 224.190 44.770 224.760 ;
        RECT 48.150 224.190 48.450 224.760 ;
        RECT 51.830 224.190 52.130 224.760 ;
        RECT 55.510 224.190 55.810 224.760 ;
        RECT 59.190 224.190 59.490 224.760 ;
        RECT 62.870 224.190 63.170 224.760 ;
        RECT 66.550 224.190 66.850 224.760 ;
        RECT 70.230 224.190 70.530 224.760 ;
        RECT 73.910 224.190 74.210 224.760 ;
        RECT 77.590 224.190 77.890 224.760 ;
        RECT 81.270 224.190 81.570 224.760 ;
        RECT 84.950 224.190 85.250 224.760 ;
        RECT 88.630 224.190 88.930 224.760 ;
        RECT 3.160 222.440 89.310 224.190 ;
        RECT 49.000 220.760 50.500 222.440 ;
        RECT 2.500 141.540 31.180 143.040 ;
        RECT 50.500 132.710 71.310 134.210 ;
        RECT 90.320 1.000 90.920 22.920 ;
        RECT 112.400 10.450 118.380 11.050 ;
        RECT 112.400 1.000 113.000 10.450 ;
        RECT 134.480 1.000 135.080 11.270 ;
        RECT 156.560 1.000 157.160 47.450 ;
  END
END tt_um_alfiero88_CurrentTrigger
END LIBRARY


magic
tech sky130A
magscale 1 2
timestamp 1716907293
<< nwell >>
rect -1949 -369 1949 369
<< pmoslvt >>
rect -1753 -150 -1613 150
rect -1555 -150 -1415 150
rect -1357 -150 -1217 150
rect -1159 -150 -1019 150
rect -961 -150 -821 150
rect -763 -150 -623 150
rect -565 -150 -425 150
rect -367 -150 -227 150
rect -169 -150 -29 150
rect 29 -150 169 150
rect 227 -150 367 150
rect 425 -150 565 150
rect 623 -150 763 150
rect 821 -150 961 150
rect 1019 -150 1159 150
rect 1217 -150 1357 150
rect 1415 -150 1555 150
rect 1613 -150 1753 150
<< pdiff >>
rect -1811 138 -1753 150
rect -1811 -138 -1799 138
rect -1765 -138 -1753 138
rect -1811 -150 -1753 -138
rect -1613 138 -1555 150
rect -1613 -138 -1601 138
rect -1567 -138 -1555 138
rect -1613 -150 -1555 -138
rect -1415 138 -1357 150
rect -1415 -138 -1403 138
rect -1369 -138 -1357 138
rect -1415 -150 -1357 -138
rect -1217 138 -1159 150
rect -1217 -138 -1205 138
rect -1171 -138 -1159 138
rect -1217 -150 -1159 -138
rect -1019 138 -961 150
rect -1019 -138 -1007 138
rect -973 -138 -961 138
rect -1019 -150 -961 -138
rect -821 138 -763 150
rect -821 -138 -809 138
rect -775 -138 -763 138
rect -821 -150 -763 -138
rect -623 138 -565 150
rect -623 -138 -611 138
rect -577 -138 -565 138
rect -623 -150 -565 -138
rect -425 138 -367 150
rect -425 -138 -413 138
rect -379 -138 -367 138
rect -425 -150 -367 -138
rect -227 138 -169 150
rect -227 -138 -215 138
rect -181 -138 -169 138
rect -227 -150 -169 -138
rect -29 138 29 150
rect -29 -138 -17 138
rect 17 -138 29 138
rect -29 -150 29 -138
rect 169 138 227 150
rect 169 -138 181 138
rect 215 -138 227 138
rect 169 -150 227 -138
rect 367 138 425 150
rect 367 -138 379 138
rect 413 -138 425 138
rect 367 -150 425 -138
rect 565 138 623 150
rect 565 -138 577 138
rect 611 -138 623 138
rect 565 -150 623 -138
rect 763 138 821 150
rect 763 -138 775 138
rect 809 -138 821 138
rect 763 -150 821 -138
rect 961 138 1019 150
rect 961 -138 973 138
rect 1007 -138 1019 138
rect 961 -150 1019 -138
rect 1159 138 1217 150
rect 1159 -138 1171 138
rect 1205 -138 1217 138
rect 1159 -150 1217 -138
rect 1357 138 1415 150
rect 1357 -138 1369 138
rect 1403 -138 1415 138
rect 1357 -150 1415 -138
rect 1555 138 1613 150
rect 1555 -138 1567 138
rect 1601 -138 1613 138
rect 1555 -150 1613 -138
rect 1753 138 1811 150
rect 1753 -138 1765 138
rect 1799 -138 1811 138
rect 1753 -150 1811 -138
<< pdiffc >>
rect -1799 -138 -1765 138
rect -1601 -138 -1567 138
rect -1403 -138 -1369 138
rect -1205 -138 -1171 138
rect -1007 -138 -973 138
rect -809 -138 -775 138
rect -611 -138 -577 138
rect -413 -138 -379 138
rect -215 -138 -181 138
rect -17 -138 17 138
rect 181 -138 215 138
rect 379 -138 413 138
rect 577 -138 611 138
rect 775 -138 809 138
rect 973 -138 1007 138
rect 1171 -138 1205 138
rect 1369 -138 1403 138
rect 1567 -138 1601 138
rect 1765 -138 1799 138
<< nsubdiff >>
rect -1913 299 -1817 333
rect 1817 299 1913 333
rect -1913 237 -1879 299
rect 1879 237 1913 299
rect -1913 -299 -1879 -237
rect 1879 -299 1913 -237
rect -1913 -333 -1817 -299
rect 1817 -333 1913 -299
<< nsubdiffcont >>
rect -1817 299 1817 333
rect -1913 -237 -1879 237
rect 1879 -237 1913 237
rect -1817 -333 1817 -299
<< poly >>
rect -1753 231 -1613 247
rect -1753 197 -1737 231
rect -1629 197 -1613 231
rect -1753 150 -1613 197
rect -1555 231 -1415 247
rect -1555 197 -1539 231
rect -1431 197 -1415 231
rect -1555 150 -1415 197
rect -1357 231 -1217 247
rect -1357 197 -1341 231
rect -1233 197 -1217 231
rect -1357 150 -1217 197
rect -1159 231 -1019 247
rect -1159 197 -1143 231
rect -1035 197 -1019 231
rect -1159 150 -1019 197
rect -961 231 -821 247
rect -961 197 -945 231
rect -837 197 -821 231
rect -961 150 -821 197
rect -763 231 -623 247
rect -763 197 -747 231
rect -639 197 -623 231
rect -763 150 -623 197
rect -565 231 -425 247
rect -565 197 -549 231
rect -441 197 -425 231
rect -565 150 -425 197
rect -367 231 -227 247
rect -367 197 -351 231
rect -243 197 -227 231
rect -367 150 -227 197
rect -169 231 -29 247
rect -169 197 -153 231
rect -45 197 -29 231
rect -169 150 -29 197
rect 29 231 169 247
rect 29 197 45 231
rect 153 197 169 231
rect 29 150 169 197
rect 227 231 367 247
rect 227 197 243 231
rect 351 197 367 231
rect 227 150 367 197
rect 425 231 565 247
rect 425 197 441 231
rect 549 197 565 231
rect 425 150 565 197
rect 623 231 763 247
rect 623 197 639 231
rect 747 197 763 231
rect 623 150 763 197
rect 821 231 961 247
rect 821 197 837 231
rect 945 197 961 231
rect 821 150 961 197
rect 1019 231 1159 247
rect 1019 197 1035 231
rect 1143 197 1159 231
rect 1019 150 1159 197
rect 1217 231 1357 247
rect 1217 197 1233 231
rect 1341 197 1357 231
rect 1217 150 1357 197
rect 1415 231 1555 247
rect 1415 197 1431 231
rect 1539 197 1555 231
rect 1415 150 1555 197
rect 1613 231 1753 247
rect 1613 197 1629 231
rect 1737 197 1753 231
rect 1613 150 1753 197
rect -1753 -197 -1613 -150
rect -1753 -231 -1737 -197
rect -1629 -231 -1613 -197
rect -1753 -247 -1613 -231
rect -1555 -197 -1415 -150
rect -1555 -231 -1539 -197
rect -1431 -231 -1415 -197
rect -1555 -247 -1415 -231
rect -1357 -197 -1217 -150
rect -1357 -231 -1341 -197
rect -1233 -231 -1217 -197
rect -1357 -247 -1217 -231
rect -1159 -197 -1019 -150
rect -1159 -231 -1143 -197
rect -1035 -231 -1019 -197
rect -1159 -247 -1019 -231
rect -961 -197 -821 -150
rect -961 -231 -945 -197
rect -837 -231 -821 -197
rect -961 -247 -821 -231
rect -763 -197 -623 -150
rect -763 -231 -747 -197
rect -639 -231 -623 -197
rect -763 -247 -623 -231
rect -565 -197 -425 -150
rect -565 -231 -549 -197
rect -441 -231 -425 -197
rect -565 -247 -425 -231
rect -367 -197 -227 -150
rect -367 -231 -351 -197
rect -243 -231 -227 -197
rect -367 -247 -227 -231
rect -169 -197 -29 -150
rect -169 -231 -153 -197
rect -45 -231 -29 -197
rect -169 -247 -29 -231
rect 29 -197 169 -150
rect 29 -231 45 -197
rect 153 -231 169 -197
rect 29 -247 169 -231
rect 227 -197 367 -150
rect 227 -231 243 -197
rect 351 -231 367 -197
rect 227 -247 367 -231
rect 425 -197 565 -150
rect 425 -231 441 -197
rect 549 -231 565 -197
rect 425 -247 565 -231
rect 623 -197 763 -150
rect 623 -231 639 -197
rect 747 -231 763 -197
rect 623 -247 763 -231
rect 821 -197 961 -150
rect 821 -231 837 -197
rect 945 -231 961 -197
rect 821 -247 961 -231
rect 1019 -197 1159 -150
rect 1019 -231 1035 -197
rect 1143 -231 1159 -197
rect 1019 -247 1159 -231
rect 1217 -197 1357 -150
rect 1217 -231 1233 -197
rect 1341 -231 1357 -197
rect 1217 -247 1357 -231
rect 1415 -197 1555 -150
rect 1415 -231 1431 -197
rect 1539 -231 1555 -197
rect 1415 -247 1555 -231
rect 1613 -197 1753 -150
rect 1613 -231 1629 -197
rect 1737 -231 1753 -197
rect 1613 -247 1753 -231
<< polycont >>
rect -1737 197 -1629 231
rect -1539 197 -1431 231
rect -1341 197 -1233 231
rect -1143 197 -1035 231
rect -945 197 -837 231
rect -747 197 -639 231
rect -549 197 -441 231
rect -351 197 -243 231
rect -153 197 -45 231
rect 45 197 153 231
rect 243 197 351 231
rect 441 197 549 231
rect 639 197 747 231
rect 837 197 945 231
rect 1035 197 1143 231
rect 1233 197 1341 231
rect 1431 197 1539 231
rect 1629 197 1737 231
rect -1737 -231 -1629 -197
rect -1539 -231 -1431 -197
rect -1341 -231 -1233 -197
rect -1143 -231 -1035 -197
rect -945 -231 -837 -197
rect -747 -231 -639 -197
rect -549 -231 -441 -197
rect -351 -231 -243 -197
rect -153 -231 -45 -197
rect 45 -231 153 -197
rect 243 -231 351 -197
rect 441 -231 549 -197
rect 639 -231 747 -197
rect 837 -231 945 -197
rect 1035 -231 1143 -197
rect 1233 -231 1341 -197
rect 1431 -231 1539 -197
rect 1629 -231 1737 -197
<< locali >>
rect -1913 299 -1817 333
rect 1817 299 1913 333
rect -1913 237 -1879 299
rect 1879 237 1913 299
rect -1753 197 -1737 231
rect -1629 197 -1613 231
rect -1555 197 -1539 231
rect -1431 197 -1415 231
rect -1357 197 -1341 231
rect -1233 197 -1217 231
rect -1159 197 -1143 231
rect -1035 197 -1019 231
rect -961 197 -945 231
rect -837 197 -821 231
rect -763 197 -747 231
rect -639 197 -623 231
rect -565 197 -549 231
rect -441 197 -425 231
rect -367 197 -351 231
rect -243 197 -227 231
rect -169 197 -153 231
rect -45 197 -29 231
rect 29 197 45 231
rect 153 197 169 231
rect 227 197 243 231
rect 351 197 367 231
rect 425 197 441 231
rect 549 197 565 231
rect 623 197 639 231
rect 747 197 763 231
rect 821 197 837 231
rect 945 197 961 231
rect 1019 197 1035 231
rect 1143 197 1159 231
rect 1217 197 1233 231
rect 1341 197 1357 231
rect 1415 197 1431 231
rect 1539 197 1555 231
rect 1613 197 1629 231
rect 1737 197 1753 231
rect -1799 138 -1765 154
rect -1799 -154 -1765 -138
rect -1601 138 -1567 154
rect -1601 -154 -1567 -138
rect -1403 138 -1369 154
rect -1403 -154 -1369 -138
rect -1205 138 -1171 154
rect -1205 -154 -1171 -138
rect -1007 138 -973 154
rect -1007 -154 -973 -138
rect -809 138 -775 154
rect -809 -154 -775 -138
rect -611 138 -577 154
rect -611 -154 -577 -138
rect -413 138 -379 154
rect -413 -154 -379 -138
rect -215 138 -181 154
rect -215 -154 -181 -138
rect -17 138 17 154
rect -17 -154 17 -138
rect 181 138 215 154
rect 181 -154 215 -138
rect 379 138 413 154
rect 379 -154 413 -138
rect 577 138 611 154
rect 577 -154 611 -138
rect 775 138 809 154
rect 775 -154 809 -138
rect 973 138 1007 154
rect 973 -154 1007 -138
rect 1171 138 1205 154
rect 1171 -154 1205 -138
rect 1369 138 1403 154
rect 1369 -154 1403 -138
rect 1567 138 1601 154
rect 1567 -154 1601 -138
rect 1765 138 1799 154
rect 1765 -154 1799 -138
rect -1753 -231 -1737 -197
rect -1629 -231 -1613 -197
rect -1555 -231 -1539 -197
rect -1431 -231 -1415 -197
rect -1357 -231 -1341 -197
rect -1233 -231 -1217 -197
rect -1159 -231 -1143 -197
rect -1035 -231 -1019 -197
rect -961 -231 -945 -197
rect -837 -231 -821 -197
rect -763 -231 -747 -197
rect -639 -231 -623 -197
rect -565 -231 -549 -197
rect -441 -231 -425 -197
rect -367 -231 -351 -197
rect -243 -231 -227 -197
rect -169 -231 -153 -197
rect -45 -231 -29 -197
rect 29 -231 45 -197
rect 153 -231 169 -197
rect 227 -231 243 -197
rect 351 -231 367 -197
rect 425 -231 441 -197
rect 549 -231 565 -197
rect 623 -231 639 -197
rect 747 -231 763 -197
rect 821 -231 837 -197
rect 945 -231 961 -197
rect 1019 -231 1035 -197
rect 1143 -231 1159 -197
rect 1217 -231 1233 -197
rect 1341 -231 1357 -197
rect 1415 -231 1431 -197
rect 1539 -231 1555 -197
rect 1613 -231 1629 -197
rect 1737 -231 1753 -197
rect -1913 -299 -1879 -237
rect 1879 -299 1913 -237
rect -1913 -333 -1817 -299
rect 1817 -333 1913 -299
<< viali >>
rect -1737 197 -1629 231
rect -1539 197 -1431 231
rect -1341 197 -1233 231
rect -1143 197 -1035 231
rect -945 197 -837 231
rect -747 197 -639 231
rect -549 197 -441 231
rect -351 197 -243 231
rect -153 197 -45 231
rect 45 197 153 231
rect 243 197 351 231
rect 441 197 549 231
rect 639 197 747 231
rect 837 197 945 231
rect 1035 197 1143 231
rect 1233 197 1341 231
rect 1431 197 1539 231
rect 1629 197 1737 231
rect -1799 -138 -1765 138
rect -1601 -138 -1567 138
rect -1403 -138 -1369 138
rect -1205 -138 -1171 138
rect -1007 -138 -973 138
rect -809 -138 -775 138
rect -611 -138 -577 138
rect -413 -138 -379 138
rect -215 -138 -181 138
rect -17 -138 17 138
rect 181 -138 215 138
rect 379 -138 413 138
rect 577 -138 611 138
rect 775 -138 809 138
rect 973 -138 1007 138
rect 1171 -138 1205 138
rect 1369 -138 1403 138
rect 1567 -138 1601 138
rect 1765 -138 1799 138
rect -1737 -231 -1629 -197
rect -1539 -231 -1431 -197
rect -1341 -231 -1233 -197
rect -1143 -231 -1035 -197
rect -945 -231 -837 -197
rect -747 -231 -639 -197
rect -549 -231 -441 -197
rect -351 -231 -243 -197
rect -153 -231 -45 -197
rect 45 -231 153 -197
rect 243 -231 351 -197
rect 441 -231 549 -197
rect 639 -231 747 -197
rect 837 -231 945 -197
rect 1035 -231 1143 -197
rect 1233 -231 1341 -197
rect 1431 -231 1539 -197
rect 1629 -231 1737 -197
<< metal1 >>
rect -1749 231 -1617 237
rect -1749 197 -1737 231
rect -1629 197 -1617 231
rect -1749 191 -1617 197
rect -1551 231 -1419 237
rect -1551 197 -1539 231
rect -1431 197 -1419 231
rect -1551 191 -1419 197
rect -1353 231 -1221 237
rect -1353 197 -1341 231
rect -1233 197 -1221 231
rect -1353 191 -1221 197
rect -1155 231 -1023 237
rect -1155 197 -1143 231
rect -1035 197 -1023 231
rect -1155 191 -1023 197
rect -957 231 -825 237
rect -957 197 -945 231
rect -837 197 -825 231
rect -957 191 -825 197
rect -759 231 -627 237
rect -759 197 -747 231
rect -639 197 -627 231
rect -759 191 -627 197
rect -561 231 -429 237
rect -561 197 -549 231
rect -441 197 -429 231
rect -561 191 -429 197
rect -363 231 -231 237
rect -363 197 -351 231
rect -243 197 -231 231
rect -363 191 -231 197
rect -165 231 -33 237
rect -165 197 -153 231
rect -45 197 -33 231
rect -165 191 -33 197
rect 33 231 165 237
rect 33 197 45 231
rect 153 197 165 231
rect 33 191 165 197
rect 231 231 363 237
rect 231 197 243 231
rect 351 197 363 231
rect 231 191 363 197
rect 429 231 561 237
rect 429 197 441 231
rect 549 197 561 231
rect 429 191 561 197
rect 627 231 759 237
rect 627 197 639 231
rect 747 197 759 231
rect 627 191 759 197
rect 825 231 957 237
rect 825 197 837 231
rect 945 197 957 231
rect 825 191 957 197
rect 1023 231 1155 237
rect 1023 197 1035 231
rect 1143 197 1155 231
rect 1023 191 1155 197
rect 1221 231 1353 237
rect 1221 197 1233 231
rect 1341 197 1353 231
rect 1221 191 1353 197
rect 1419 231 1551 237
rect 1419 197 1431 231
rect 1539 197 1551 231
rect 1419 191 1551 197
rect 1617 231 1749 237
rect 1617 197 1629 231
rect 1737 197 1749 231
rect 1617 191 1749 197
rect -1805 138 -1759 150
rect -1805 -138 -1799 138
rect -1765 -138 -1759 138
rect -1805 -150 -1759 -138
rect -1607 138 -1561 150
rect -1607 -138 -1601 138
rect -1567 -138 -1561 138
rect -1607 -150 -1561 -138
rect -1409 138 -1363 150
rect -1409 -138 -1403 138
rect -1369 -138 -1363 138
rect -1409 -150 -1363 -138
rect -1211 138 -1165 150
rect -1211 -138 -1205 138
rect -1171 -138 -1165 138
rect -1211 -150 -1165 -138
rect -1013 138 -967 150
rect -1013 -138 -1007 138
rect -973 -138 -967 138
rect -1013 -150 -967 -138
rect -815 138 -769 150
rect -815 -138 -809 138
rect -775 -138 -769 138
rect -815 -150 -769 -138
rect -617 138 -571 150
rect -617 -138 -611 138
rect -577 -138 -571 138
rect -617 -150 -571 -138
rect -419 138 -373 150
rect -419 -138 -413 138
rect -379 -138 -373 138
rect -419 -150 -373 -138
rect -221 138 -175 150
rect -221 -138 -215 138
rect -181 -138 -175 138
rect -221 -150 -175 -138
rect -23 138 23 150
rect -23 -138 -17 138
rect 17 -138 23 138
rect -23 -150 23 -138
rect 175 138 221 150
rect 175 -138 181 138
rect 215 -138 221 138
rect 175 -150 221 -138
rect 373 138 419 150
rect 373 -138 379 138
rect 413 -138 419 138
rect 373 -150 419 -138
rect 571 138 617 150
rect 571 -138 577 138
rect 611 -138 617 138
rect 571 -150 617 -138
rect 769 138 815 150
rect 769 -138 775 138
rect 809 -138 815 138
rect 769 -150 815 -138
rect 967 138 1013 150
rect 967 -138 973 138
rect 1007 -138 1013 138
rect 967 -150 1013 -138
rect 1165 138 1211 150
rect 1165 -138 1171 138
rect 1205 -138 1211 138
rect 1165 -150 1211 -138
rect 1363 138 1409 150
rect 1363 -138 1369 138
rect 1403 -138 1409 138
rect 1363 -150 1409 -138
rect 1561 138 1607 150
rect 1561 -138 1567 138
rect 1601 -138 1607 138
rect 1561 -150 1607 -138
rect 1759 138 1805 150
rect 1759 -138 1765 138
rect 1799 -138 1805 138
rect 1759 -150 1805 -138
rect -1749 -197 -1617 -191
rect -1749 -231 -1737 -197
rect -1629 -231 -1617 -197
rect -1749 -237 -1617 -231
rect -1551 -197 -1419 -191
rect -1551 -231 -1539 -197
rect -1431 -231 -1419 -197
rect -1551 -237 -1419 -231
rect -1353 -197 -1221 -191
rect -1353 -231 -1341 -197
rect -1233 -231 -1221 -197
rect -1353 -237 -1221 -231
rect -1155 -197 -1023 -191
rect -1155 -231 -1143 -197
rect -1035 -231 -1023 -197
rect -1155 -237 -1023 -231
rect -957 -197 -825 -191
rect -957 -231 -945 -197
rect -837 -231 -825 -197
rect -957 -237 -825 -231
rect -759 -197 -627 -191
rect -759 -231 -747 -197
rect -639 -231 -627 -197
rect -759 -237 -627 -231
rect -561 -197 -429 -191
rect -561 -231 -549 -197
rect -441 -231 -429 -197
rect -561 -237 -429 -231
rect -363 -197 -231 -191
rect -363 -231 -351 -197
rect -243 -231 -231 -197
rect -363 -237 -231 -231
rect -165 -197 -33 -191
rect -165 -231 -153 -197
rect -45 -231 -33 -197
rect -165 -237 -33 -231
rect 33 -197 165 -191
rect 33 -231 45 -197
rect 153 -231 165 -197
rect 33 -237 165 -231
rect 231 -197 363 -191
rect 231 -231 243 -197
rect 351 -231 363 -197
rect 231 -237 363 -231
rect 429 -197 561 -191
rect 429 -231 441 -197
rect 549 -231 561 -197
rect 429 -237 561 -231
rect 627 -197 759 -191
rect 627 -231 639 -197
rect 747 -231 759 -197
rect 627 -237 759 -231
rect 825 -197 957 -191
rect 825 -231 837 -197
rect 945 -231 957 -197
rect 825 -237 957 -231
rect 1023 -197 1155 -191
rect 1023 -231 1035 -197
rect 1143 -231 1155 -197
rect 1023 -237 1155 -231
rect 1221 -197 1353 -191
rect 1221 -231 1233 -197
rect 1341 -231 1353 -197
rect 1221 -237 1353 -231
rect 1419 -197 1551 -191
rect 1419 -231 1431 -197
rect 1539 -231 1551 -197
rect 1419 -237 1551 -231
rect 1617 -197 1749 -191
rect 1617 -231 1629 -197
rect 1737 -231 1749 -197
rect 1617 -237 1749 -231
<< properties >>
string FIXED_BBOX -1896 -316 1896 316
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1.5 l 0.7 m 1 nf 18 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1716974663
<< error_s >>
rect 10936 6462 10998 6468
rect 11064 6462 11126 6468
rect 11192 6462 11254 6468
rect 11320 6462 11382 6468
rect 11448 6462 11510 6468
rect 11576 6462 11638 6468
rect 11704 6462 11766 6468
rect 10936 6428 10948 6462
rect 11064 6428 11076 6462
rect 11192 6428 11204 6462
rect 11320 6428 11332 6462
rect 11448 6428 11460 6462
rect 11576 6428 11588 6462
rect 11704 6428 11716 6462
rect 10936 6422 10998 6428
rect 11064 6422 11126 6428
rect 11192 6422 11254 6428
rect 11320 6422 11382 6428
rect 11448 6422 11510 6428
rect 11576 6422 11638 6428
rect 11704 6422 11766 6428
rect 13378 6348 13440 6354
rect 13506 6348 13568 6354
rect 13634 6348 13696 6354
rect 13378 6314 13390 6348
rect 13506 6314 13518 6348
rect 13634 6314 13646 6348
rect 13378 6308 13440 6314
rect 13506 6308 13568 6314
rect 13634 6308 13696 6314
rect 19982 5934 20044 5940
rect 20110 5934 20172 5940
rect 20238 5934 20300 5940
rect 20366 5934 20428 5940
rect 20494 5934 20556 5940
rect 20622 5934 20684 5940
rect 10936 5906 10998 5912
rect 11064 5906 11126 5912
rect 11192 5906 11254 5912
rect 11320 5906 11382 5912
rect 11448 5906 11510 5912
rect 11576 5906 11638 5912
rect 11704 5906 11766 5912
rect 10936 5872 10948 5906
rect 11064 5872 11076 5906
rect 11192 5872 11204 5906
rect 11320 5872 11332 5906
rect 11448 5872 11460 5906
rect 11576 5872 11588 5906
rect 11704 5872 11716 5906
rect 19982 5900 19994 5934
rect 20110 5900 20122 5934
rect 20238 5900 20250 5934
rect 20366 5900 20378 5934
rect 20494 5900 20506 5934
rect 20622 5900 20634 5934
rect 19982 5894 20044 5900
rect 20110 5894 20172 5900
rect 20238 5894 20300 5900
rect 20366 5894 20428 5900
rect 20494 5894 20556 5900
rect 20622 5894 20684 5900
rect 13378 5886 13440 5892
rect 13506 5886 13568 5892
rect 13634 5886 13696 5892
rect 10936 5866 10998 5872
rect 11064 5866 11126 5872
rect 11192 5866 11254 5872
rect 11320 5866 11382 5872
rect 11448 5866 11510 5872
rect 11576 5866 11638 5872
rect 11704 5866 11766 5872
rect 13378 5852 13390 5886
rect 13506 5852 13518 5886
rect 13634 5852 13646 5886
rect 13378 5846 13440 5852
rect 13506 5846 13568 5852
rect 13634 5846 13696 5852
rect 17200 5734 17262 5740
rect 18474 5734 18536 5740
rect 18602 5734 18664 5740
rect 18730 5734 18792 5740
rect 17200 5700 17212 5734
rect 18474 5700 18486 5734
rect 18602 5700 18614 5734
rect 18730 5700 18742 5734
rect 17200 5694 17262 5700
rect 18474 5694 18536 5700
rect 18602 5694 18664 5700
rect 18730 5694 18792 5700
rect 17200 5206 17262 5212
rect 18474 5206 18536 5212
rect 18602 5206 18664 5212
rect 18730 5206 18792 5212
rect 19982 5206 20044 5212
rect 20110 5206 20172 5212
rect 20238 5206 20300 5212
rect 20366 5206 20428 5212
rect 20494 5206 20556 5212
rect 20622 5206 20684 5212
rect 17200 5172 17212 5206
rect 18474 5172 18486 5206
rect 18602 5172 18614 5206
rect 18730 5172 18742 5206
rect 19982 5172 19994 5206
rect 20110 5172 20122 5206
rect 20238 5172 20250 5206
rect 20366 5196 20378 5206
rect 20494 5172 20506 5206
rect 20622 5172 20634 5206
rect 17200 5166 17262 5172
rect 18474 5166 18536 5172
rect 18602 5166 18664 5172
rect 18730 5166 18792 5172
rect 19982 5166 20044 5172
rect 20110 5166 20172 5172
rect 20238 5166 20252 5172
rect 20494 5166 20556 5172
rect 20622 5166 20684 5172
rect 20106 3664 20164 3670
rect 20106 3630 20118 3664
rect 20106 3624 20164 3630
rect 18556 3386 18614 3392
rect 18556 3352 18568 3386
rect 18556 3346 18614 3352
rect 17162 3286 17220 3292
rect 17162 3252 17174 3286
rect 17162 3246 17220 3252
rect 17162 2976 17220 2982
rect 18460 2976 18518 2982
rect 17162 2942 17174 2976
rect 18460 2942 18472 2976
rect 20010 2954 20068 2960
rect 20202 2954 20260 2960
rect 17162 2936 17220 2942
rect 18460 2936 18518 2942
rect 20010 2920 20022 2954
rect 20202 2920 20214 2954
rect 20010 2914 20068 2920
rect 20202 2914 20260 2920
<< error_ps >>
rect 20366 5172 20378 5196
rect 20252 5166 20300 5172
rect 20366 5166 20428 5172
<< viali >>
rect 246 9102 982 9142
rect 126 6584 166 7364
rect 4010 7212 7630 7272
rect 122 4756 166 5526
rect 3256 2836 5312 2884
rect 222 2726 960 2768
<< metal1 >>
rect -812 9296 21028 10100
rect -812 8898 -340 9296
rect 154 9142 1078 9296
rect 154 9102 246 9142
rect 982 9102 1078 9142
rect 154 9096 1078 9102
rect 1275 9038 1385 9039
rect 302 8988 1385 9038
rect -812 8392 302 8898
rect 1240 8812 1385 8988
rect 922 8582 1385 8812
rect -812 7372 -340 8392
rect 1240 8308 1385 8582
rect 302 8258 1385 8308
rect 1275 7949 1385 8258
rect 1275 7839 1531 7949
rect 1422 7772 1530 7839
rect 1416 7664 1422 7772
rect 1530 7664 1536 7772
rect 2980 7590 3624 9296
rect -812 7364 180 7372
rect 1592 7368 1654 7369
rect -812 6584 126 7364
rect 166 6584 180 7364
rect 280 7306 1654 7368
rect 352 7170 362 7266
rect 418 7170 428 7266
rect 610 7170 620 7266
rect 676 7170 686 7266
rect 864 7170 874 7266
rect 930 7170 940 7266
rect 1120 7170 1130 7266
rect 1186 7170 1196 7266
rect 1414 6796 1530 6802
rect 1592 6796 1654 7306
rect 2979 7272 7642 7590
rect 3984 7212 4010 7272
rect 7630 7212 7642 7272
rect 3984 7198 7642 7212
rect 4052 7104 8098 7168
rect 3988 6964 3998 7070
rect 4056 6964 4066 7070
rect 4384 6964 4394 7070
rect 4452 6964 4462 7070
rect 4780 6964 4790 7070
rect 4848 6964 4858 7070
rect 5174 6964 5184 7070
rect 5242 6964 5252 7070
rect 5570 6964 5580 7070
rect 5638 6964 5648 7070
rect 5968 6964 5978 7070
rect 6036 6964 6046 7070
rect 6364 6964 6374 7070
rect 6432 6964 6442 7070
rect 6758 6964 6768 7070
rect 6826 6964 6836 7070
rect 7156 6964 7166 7070
rect 7224 6964 7234 7070
rect 7552 6964 7562 7070
rect 7620 6964 7630 7070
rect 238 6690 248 6786
rect 304 6690 314 6786
rect 482 6686 492 6782
rect 548 6686 558 6782
rect 736 6686 746 6782
rect 802 6686 812 6782
rect 994 6686 1004 6782
rect 1060 6686 1070 6782
rect 1530 6680 1654 6796
rect 4186 6772 4196 6878
rect 4254 6772 4264 6878
rect 4580 6772 4590 6878
rect 4648 6772 4658 6878
rect 4976 6772 4986 6878
rect 5044 6772 5054 6878
rect 5374 6772 5384 6878
rect 5442 6772 5452 6878
rect 5770 6772 5780 6878
rect 5838 6772 5848 6878
rect 6164 6772 6174 6878
rect 6232 6772 6242 6878
rect 6560 6772 6570 6878
rect 6628 6772 6638 6878
rect 6956 6772 6966 6878
rect 7024 6772 7034 6878
rect 7352 6772 7362 6878
rect 7420 6772 7430 6878
rect 8026 6726 8090 7104
rect 21630 6864 21830 7064
rect 1414 6664 1654 6680
rect 1414 6636 1658 6664
rect 4056 6662 8102 6726
rect -812 6570 180 6584
rect 280 6574 1658 6636
rect -354 6568 180 6570
rect -854 5926 677 6239
rect 990 5926 996 6239
rect -326 5582 172 5584
rect -782 5526 172 5582
rect 1538 5538 1658 6574
rect 8026 5594 8090 6662
rect -782 4756 122 5526
rect 166 4756 172 5526
rect 366 5468 1658 5538
rect 4044 5530 8090 5594
rect 228 5342 238 5440
rect 296 5342 306 5440
rect 416 5342 426 5440
rect 484 5342 494 5440
rect 608 5342 618 5440
rect 676 5342 686 5440
rect 800 5342 810 5440
rect 868 5342 878 5440
rect 1538 5293 1658 5468
rect 1158 5179 1164 5293
rect 1278 5179 1658 5293
rect 320 4854 330 4952
rect 388 4854 398 4952
rect 512 4854 522 4952
rect 580 4854 590 4952
rect 704 4854 714 4952
rect 772 4854 782 4952
rect 896 4854 906 4952
rect 964 4854 974 4952
rect 1538 4808 1658 5179
rect 8026 5162 8090 5530
rect 4044 5098 8090 5162
rect -782 4718 172 4756
rect 276 4738 1658 4808
rect 1538 4736 1658 4738
rect -782 3502 -310 4718
rect 1176 4386 1288 4392
rect 1288 4382 1650 4386
rect 1288 4274 1666 4382
rect 9188 4274 9388 4474
rect 21720 4300 21920 4500
rect 1176 4268 1288 4274
rect 1530 3922 1666 4274
rect 2570 3922 5284 3924
rect 1530 3856 5284 3922
rect 1530 3736 2638 3856
rect 1530 3598 1666 3736
rect 290 3538 1666 3598
rect -782 2916 284 3502
rect 894 3220 978 3502
rect 894 3219 1144 3220
rect 1530 3219 1666 3538
rect 894 3053 1666 3219
rect 894 3052 1144 3053
rect 894 2922 978 3052
rect -782 2486 -310 2916
rect 1530 2878 1666 3053
rect 2570 2996 2638 3736
rect 3256 3684 3266 3810
rect 3330 3684 3340 3810
rect 4572 3684 4582 3810
rect 4646 3684 4656 3810
rect 3910 3038 3920 3164
rect 3984 3038 3994 3164
rect 5232 3038 5242 3164
rect 5306 3038 5316 3164
rect 2570 2946 5244 2996
rect 292 2830 1666 2878
rect 3244 2884 5332 2890
rect 3244 2836 3256 2884
rect 5312 2836 5332 2884
rect 170 2768 1018 2774
rect 170 2726 222 2768
rect 960 2726 1018 2768
rect 170 2486 1018 2726
rect 3244 2486 5332 2836
rect -784 1682 21056 2486
<< via1 >>
rect 1422 7664 1530 7772
rect 362 7170 418 7266
rect 620 7170 676 7266
rect 874 7170 930 7266
rect 1130 7170 1186 7266
rect 3998 6964 4056 7070
rect 4394 6964 4452 7070
rect 4790 6964 4848 7070
rect 5184 6964 5242 7070
rect 5580 6964 5638 7070
rect 5978 6964 6036 7070
rect 6374 6964 6432 7070
rect 6768 6964 6826 7070
rect 7166 6964 7224 7070
rect 7562 6964 7620 7070
rect 248 6690 304 6786
rect 492 6686 548 6782
rect 746 6686 802 6782
rect 1004 6686 1060 6782
rect 1414 6680 1530 6796
rect 4196 6772 4254 6878
rect 4590 6772 4648 6878
rect 4986 6772 5044 6878
rect 5384 6772 5442 6878
rect 5780 6772 5838 6878
rect 6174 6772 6232 6878
rect 6570 6772 6628 6878
rect 6966 6772 7024 6878
rect 7362 6772 7420 6878
rect 677 5926 990 6239
rect 238 5342 296 5440
rect 426 5342 484 5440
rect 618 5342 676 5440
rect 810 5342 868 5440
rect 1164 5179 1278 5293
rect 330 4854 388 4952
rect 522 4854 580 4952
rect 714 4854 772 4952
rect 906 4854 964 4952
rect 1176 4274 1288 4386
rect 3266 3684 3330 3810
rect 4582 3684 4646 3810
rect 3920 3038 3984 3164
rect 5242 3038 5306 3164
<< metal2 >>
rect 1422 7772 1530 7778
rect 362 7272 418 7276
rect 620 7272 676 7276
rect 874 7272 930 7276
rect 1130 7272 1186 7276
rect 1422 7272 1530 7664
rect 350 7266 1530 7272
rect 350 7170 362 7266
rect 418 7170 620 7266
rect 676 7170 874 7266
rect 930 7170 1130 7266
rect 1186 7170 1530 7266
rect 350 7164 1530 7170
rect 362 7160 418 7164
rect 620 7160 676 7164
rect 874 7160 930 7164
rect 1130 7160 1186 7164
rect 2519 7078 3262 7168
rect 3998 7078 4056 7080
rect 4394 7078 4452 7080
rect 4790 7078 4848 7080
rect 5184 7078 5242 7080
rect 5580 7078 5638 7080
rect 5978 7078 6036 7080
rect 6374 7078 6432 7080
rect 6768 7078 6826 7080
rect 7166 7078 7224 7080
rect 7562 7078 7620 7080
rect 2519 7070 7627 7078
rect 2519 6964 3998 7070
rect 4056 6964 4394 7070
rect 4452 6964 4790 7070
rect 4848 6964 5184 7070
rect 5242 6964 5580 7070
rect 5638 6964 5978 7070
rect 6036 6964 6374 7070
rect 6432 6964 6768 7070
rect 6826 6964 7166 7070
rect 7224 6964 7562 7070
rect 7620 6964 7627 7070
rect 2519 6944 7627 6964
rect 2519 6855 3262 6944
rect 4196 6878 4254 6888
rect 246 6786 1414 6796
rect 246 6690 248 6786
rect 304 6782 1414 6786
rect 304 6690 492 6782
rect 246 6686 492 6690
rect 548 6686 746 6782
rect 802 6686 1004 6782
rect 1060 6686 1414 6782
rect 246 6680 1414 6686
rect 1530 6680 1536 6796
rect 492 6676 548 6680
rect 746 6676 802 6680
rect 1004 6676 1060 6680
rect 677 6239 990 6245
rect 2519 6239 2832 6855
rect 4196 6762 4254 6772
rect 4590 6878 4648 6888
rect 4590 6762 4648 6772
rect 4986 6878 5044 6888
rect 4986 6762 5044 6772
rect 5384 6878 5442 6888
rect 5384 6762 5442 6772
rect 5780 6878 5838 6888
rect 5780 6762 5838 6772
rect 6174 6878 6232 6888
rect 6174 6762 6232 6772
rect 6570 6878 6628 6888
rect 6570 6762 6628 6772
rect 6966 6878 7024 6888
rect 6966 6762 7024 6772
rect 7362 6878 7420 6888
rect 7362 6762 7420 6772
rect 990 5926 2832 6239
rect 677 5920 990 5926
rect 238 5440 1278 5450
rect 296 5342 426 5440
rect 484 5342 618 5440
rect 676 5342 810 5440
rect 868 5342 1278 5440
rect 238 5336 1278 5342
rect 238 5332 296 5336
rect 426 5332 484 5336
rect 618 5332 676 5336
rect 810 5332 868 5336
rect 1164 5293 1278 5336
rect 1164 5173 1278 5179
rect 330 4952 1288 4962
rect 388 4854 522 4952
rect 580 4854 714 4952
rect 772 4854 906 4952
rect 964 4854 1288 4952
rect 330 4850 1288 4854
rect 330 4844 388 4850
rect 522 4844 580 4850
rect 714 4844 772 4850
rect 906 4844 964 4850
rect 1176 4386 1288 4850
rect 1170 4274 1176 4386
rect 1288 4274 1294 4386
rect 3266 3810 3330 3820
rect 3266 3674 3330 3684
rect 4582 3810 4646 3820
rect 4582 3674 4646 3684
rect 3920 3164 3984 3174
rect 3920 3028 3984 3038
rect 5242 3164 5306 3174
rect 5242 3028 5306 3038
use sky130_fd_pr__nfet_01v8_lvt_BSZA4P  XM1
timestamp 1716907293
transform 1 0 18404 0 1 6978
box -554 -310 554 310
use sky130_fd_pr__nfet_01v8_lvt_BSZA4P  XM2
timestamp 1716907293
transform 1 0 12398 0 1 3008
box -554 -310 554 310
use sky130_fd_pr__pfet_01v8_lvt_366EDY  XM3
timestamp 1716907293
transform 1 0 11351 0 1 6167
box -615 -433 615 433
use sky130_fd_pr__pfet_01v8_lvt_ET6TZU  XM4
timestamp 1716907293
transform 1 0 5809 0 1 5349
box -1949 -369 1949 369
use sky130_fd_pr__pfet_01v8_lvt_ET6TZU  XM5
timestamp 1716907293
transform 1 0 5809 0 1 6915
box -1949 -369 1949 369
use sky130_fd_pr__pfet_01v8_lvt_CE5TV5  XM6
timestamp 1716907293
transform 1 0 7662 0 1 8533
box -3128 -419 3128 419
use sky130_fd_pr__pfet_01v8_lvt_QBWM73  XM7
timestamp 1716907293
transform 1 0 13537 0 1 6100
box -359 -386 359 386
use sky130_fd_pr__nfet_01v8_lvt_XWWVRJ  XM8
timestamp 1716907293
transform 1 0 12418 0 1 4430
box -854 -310 854 310
use sky130_fd_pr__pfet_01v8_lvt_CEZKS5  XM9
timestamp 1716907293
transform 1 0 18695 0 1 8553
box -2141 -419 2141 419
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XM10
timestamp 1716907293
transform 1 0 17191 0 1 3114
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_lvt_4QFWD3  XM11
timestamp 1716907293
transform 1 0 17231 0 1 5453
box -231 -419 231 419
use sky130_fd_pr__pfet_01v8_lvt_4QPJD3  XM12
timestamp 1716907293
transform 1 0 18633 0 1 5453
box -359 -419 359 419
use sky130_fd_pr__nfet_01v8_lvt_CW7PBK  XM13
timestamp 1716907293
transform 1 0 18537 0 1 3164
box -263 -360 263 360
use sky130_fd_pr__pfet_01v8_lvt_4QK4B3  XM14
timestamp 1716907293
transform 1 0 20333 0 1 5553
box -551 -519 551 519
use sky130_fd_pr__nfet_01v8_lvt_E5PS5K  XM15
timestamp 1716907293
transform 1 0 20135 0 1 3292
box -311 -510 311 510
use sky130_fd_pr__nfet_01v8_lvt_HEVHEL  XM16
timestamp 1716907293
transform 1 0 7404 0 1 3436
box -1154 -610 1154 610
use sky130_fd_pr__nfet_01v8_lvt_HEVHEL  XM17
timestamp 1716907293
transform 1 0 4284 0 1 3424
box -1154 -610 1154 610
use sky130_fd_pr__nfet_01v8_lvt_UJF2WX  XM18
timestamp 1716907293
transform 1 0 592 0 1 3208
box -496 -510 496 510
use sky130_fd_pr__pfet_01v8_lvt_CEYSV5  XM19
timestamp 1716907293
transform 1 0 614 0 1 8653
box -496 -519 496 519
use sky130_fd_pr__nfet_01v8_lvt_95PS5T  XM20
timestamp 1716907293
transform 1 0 599 0 1 5140
box -503 -510 503 510
use sky130_fd_pr__pfet_01v8_lvt_4QPHR2  XM21
timestamp 1716907293
transform 1 0 711 0 1 6975
box -615 -519 615 519
<< labels >>
flabel metal1 -704 1944 -504 2144 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 21720 4300 21920 4500 0 FreeSans 256 0 0 0 out
port 4 nsew
flabel metal1 21630 6864 21830 7064 0 FreeSans 256 0 0 0 in
port 5 nsew
flabel metal1 9188 4274 9388 4474 0 FreeSans 256 0 0 0 vgf
port 3 nsew
flabel metal1 -798 5982 -598 6182 0 FreeSans 256 0 0 0 vref
port 2 nsew
flabel metal1 -686 9592 -486 9792 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 1530 3736 2638 3922 0 FreeSans 1600 0 0 0 i_n
flabel metal1 1538 4736 1658 6664 0 FreeSans 1600 0 0 0 dcon
<< end >>

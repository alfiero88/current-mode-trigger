magic
tech sky130A
timestamp 1716907293
<< pwell >>
rect -577 -305 577 305
<< nmoslvt >>
rect -479 -200 -179 200
rect -150 -200 150 200
rect 179 -200 479 200
<< ndiff >>
rect -508 194 -479 200
rect -508 -194 -502 194
rect -485 -194 -479 194
rect -508 -200 -479 -194
rect -179 194 -150 200
rect -179 -194 -173 194
rect -156 -194 -150 194
rect -179 -200 -150 -194
rect 150 194 179 200
rect 150 -194 156 194
rect 173 -194 179 194
rect 150 -200 179 -194
rect 479 194 508 200
rect 479 -194 485 194
rect 502 -194 508 194
rect 479 -200 508 -194
<< ndiffc >>
rect -502 -194 -485 194
rect -173 -194 -156 194
rect 156 -194 173 194
rect 485 -194 502 194
<< psubdiff >>
rect -559 270 -511 287
rect 511 270 559 287
rect -559 239 -542 270
rect 542 239 559 270
rect -559 -270 -542 -239
rect 542 -270 559 -239
rect -559 -287 -511 -270
rect 511 -287 559 -270
<< psubdiffcont >>
rect -511 270 511 287
rect -559 -239 -542 239
rect 542 -239 559 239
rect -511 -287 511 -270
<< poly >>
rect -479 236 -179 244
rect -479 219 -471 236
rect -187 219 -179 236
rect -479 200 -179 219
rect -150 236 150 244
rect -150 219 -142 236
rect 142 219 150 236
rect -150 200 150 219
rect 179 236 479 244
rect 179 219 187 236
rect 471 219 479 236
rect 179 200 479 219
rect -479 -219 -179 -200
rect -479 -236 -471 -219
rect -187 -236 -179 -219
rect -479 -244 -179 -236
rect -150 -219 150 -200
rect -150 -236 -142 -219
rect 142 -236 150 -219
rect -150 -244 150 -236
rect 179 -219 479 -200
rect 179 -236 187 -219
rect 471 -236 479 -219
rect 179 -244 479 -236
<< polycont >>
rect -471 219 -187 236
rect -142 219 142 236
rect 187 219 471 236
rect -471 -236 -187 -219
rect -142 -236 142 -219
rect 187 -236 471 -219
<< locali >>
rect -559 270 -511 287
rect 511 270 559 287
rect -559 239 -542 270
rect 542 239 559 270
rect -479 219 -471 236
rect -187 219 -179 236
rect -150 219 -142 236
rect 142 219 150 236
rect 179 219 187 236
rect 471 219 479 236
rect -502 194 -485 202
rect -502 -202 -485 -194
rect -173 194 -156 202
rect -173 -202 -156 -194
rect 156 194 173 202
rect 156 -202 173 -194
rect 485 194 502 202
rect 485 -202 502 -194
rect -479 -236 -471 -219
rect -187 -236 -179 -219
rect -150 -236 -142 -219
rect 142 -236 150 -219
rect 179 -236 187 -219
rect 471 -236 479 -219
rect -559 -270 -542 -239
rect 542 -270 559 -239
rect -559 -287 -511 -270
rect 511 -287 559 -270
<< viali >>
rect -471 219 -187 236
rect -142 219 142 236
rect 187 219 471 236
rect -502 -194 -485 194
rect -173 -194 -156 194
rect 156 -194 173 194
rect 485 -194 502 194
rect -471 -236 -187 -219
rect -142 -236 142 -219
rect 187 -236 471 -219
<< metal1 >>
rect -477 236 -181 239
rect -477 219 -471 236
rect -187 219 -181 236
rect -477 216 -181 219
rect -148 236 148 239
rect -148 219 -142 236
rect 142 219 148 236
rect -148 216 148 219
rect 181 236 477 239
rect 181 219 187 236
rect 471 219 477 236
rect 181 216 477 219
rect -505 194 -482 200
rect -505 -194 -502 194
rect -485 -194 -482 194
rect -505 -200 -482 -194
rect -176 194 -153 200
rect -176 -194 -173 194
rect -156 -194 -153 194
rect -176 -200 -153 -194
rect 153 194 176 200
rect 153 -194 156 194
rect 173 -194 176 194
rect 153 -200 176 -194
rect 482 194 505 200
rect 482 -194 485 194
rect 502 -194 505 194
rect 482 -200 505 -194
rect -477 -219 -181 -216
rect -477 -236 -471 -219
rect -187 -236 -181 -219
rect -477 -239 -181 -236
rect -148 -219 148 -216
rect -148 -236 -142 -219
rect 142 -236 148 -219
rect -148 -239 148 -236
rect 181 -219 477 -216
rect 181 -236 187 -219
rect 471 -236 477 -219
rect 181 -239 477 -236
<< properties >>
string FIXED_BBOX -550 -278 550 278
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 4.0 l 3.0 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

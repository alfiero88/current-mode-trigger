magic
tech sky130A
magscale 1 2
timestamp 1717087242
<< metal1 >>
rect 25804 32445 26395 32472
rect 25804 31908 25831 32445
rect 26368 31908 26395 32445
rect 18142 30691 18771 30735
rect 17497 30616 18771 30691
rect 17497 30224 17572 30616
rect 17964 30224 18771 30616
rect 17497 30149 18771 30224
rect 18142 27976 18771 30149
rect 23784 29498 24060 29504
rect 22386 29222 23784 29498
rect 22386 28212 22662 29222
rect 23784 29216 24060 29222
rect 25804 27995 26395 31908
rect 19344 16587 19659 16593
rect 19659 16272 20457 16587
rect 19344 16266 19659 16272
rect 23630 9745 23923 10510
rect 23624 9452 23630 9745
rect 23923 9452 23929 9745
rect 21609 7717 21932 9031
rect 21603 7394 21609 7717
rect 21932 7394 21938 7717
<< via1 >>
rect 25831 31908 26368 32445
rect 17572 30224 17964 30616
rect 23784 29222 24060 29498
rect 19344 16272 19659 16587
rect 23630 9452 23923 9745
rect 21609 7394 21932 7717
<< metal2 >>
rect 25831 32445 26368 32451
rect 15845 32352 16182 32354
rect 17499 32352 25831 32445
rect 15838 32345 25831 32352
rect 15838 32008 15845 32345
rect 16182 32008 25831 32345
rect 15838 32001 25831 32008
rect 15845 31999 16182 32001
rect 17499 31908 25831 32001
rect 25831 31902 26368 31908
rect 15179 30570 15469 30574
rect 16632 30570 17572 30616
rect 15174 30565 17572 30570
rect 15174 30275 15179 30565
rect 15469 30275 17572 30565
rect 15174 30270 17572 30275
rect 15179 30266 15469 30270
rect 16632 30224 17572 30270
rect 17964 30224 17970 30616
rect 24265 29498 24531 29502
rect 23778 29222 23784 29498
rect 24060 29493 24536 29498
rect 24060 29227 24265 29493
rect 24531 29227 24536 29493
rect 24060 29222 24536 29227
rect 24265 29218 24531 29222
rect 15047 16272 19344 16587
rect 19659 16272 19665 16587
rect 15047 13510 15362 16272
rect 15043 13205 15052 13510
rect 15357 13205 15366 13510
rect 15047 13200 15362 13205
rect 23630 9745 23923 9751
rect 23630 7765 23923 9452
rect 21609 7717 21932 7723
rect 23626 7482 23635 7765
rect 23918 7482 23927 7765
rect 23630 7477 23923 7482
rect 21609 6644 21932 7394
rect 21605 6331 21614 6644
rect 21927 6331 21936 6644
rect 21609 6326 21932 6331
<< via2 >>
rect 15845 32008 16182 32345
rect 15179 30275 15469 30565
rect 24265 29227 24531 29493
rect 15052 13205 15357 13510
rect 23635 7482 23918 7765
rect 21614 6331 21927 6644
<< metal3 >>
rect 14963 32345 16187 32350
rect 6091 32326 6389 32331
rect 14963 32326 15845 32345
rect 6090 32325 15845 32326
rect 6090 32027 6091 32325
rect 6389 32027 15845 32325
rect 6090 32026 15845 32027
rect 6091 32021 6389 32026
rect 14963 32008 15845 32026
rect 16182 32008 16187 32345
rect 14963 32003 16187 32008
rect 14235 30570 14533 30575
rect 14234 30569 15474 30570
rect 14234 30271 14235 30569
rect 14533 30565 15474 30569
rect 14533 30275 15179 30565
rect 15469 30275 15474 30565
rect 14533 30271 15474 30275
rect 14234 30270 15474 30271
rect 14235 30265 14533 30270
rect 24767 29498 25041 29503
rect 24260 29497 25042 29498
rect 24260 29493 24767 29497
rect 24260 29227 24265 29493
rect 24531 29227 24767 29493
rect 24260 29223 24767 29227
rect 25041 29223 25042 29497
rect 24260 29222 25042 29223
rect 24767 29217 25041 29222
rect 15047 13510 15362 13515
rect 15047 13205 15052 13510
rect 15357 13205 15362 13510
rect 15047 11920 15362 13205
rect 15042 11607 15048 11920
rect 15361 11607 15367 11920
rect 15047 11606 15362 11607
rect 23630 7765 23923 7770
rect 23630 7482 23635 7765
rect 23918 7482 23923 7765
rect 23630 6735 23923 7482
rect 21609 6644 21932 6649
rect 21609 6331 21614 6644
rect 21927 6331 21932 6644
rect 23625 6444 23631 6735
rect 23922 6444 23928 6735
rect 23630 6443 23923 6444
rect 21609 5608 21932 6331
rect 21604 5287 21610 5608
rect 21931 5287 21937 5608
rect 21609 5286 21932 5287
<< via3 >>
rect 6091 32027 6389 32325
rect 14235 30271 14533 30569
rect 24767 29223 25041 29497
rect 15048 11607 15361 11920
rect 23631 6444 23922 6735
rect 21610 5287 21931 5608
<< metal4 >>
rect 798 44714 858 45152
rect 1534 44714 1594 45152
rect 2270 44714 2330 45152
rect 3006 44714 3066 45152
rect 3742 44714 3802 45152
rect 4478 44714 4538 45152
rect 5214 44714 5274 45152
rect 5950 44714 6010 45152
rect 6686 44714 6746 45152
rect 7422 44714 7482 45152
rect 8158 44714 8218 45152
rect 8894 44714 8954 45152
rect 9630 44714 9690 45152
rect 10366 44714 10426 45152
rect 11102 44714 11162 45152
rect 11838 44714 11898 45152
rect 12574 44714 12634 45152
rect 13310 44714 13370 45152
rect 14046 44714 14106 45152
rect 14782 44714 14842 45152
rect 15518 44714 15578 45152
rect 16254 44714 16314 45152
rect 16990 44714 17050 45152
rect 17726 44714 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 752 44430 17788 44714
rect 200 32326 500 44152
rect 200 32325 6390 32326
rect 200 32027 6091 32325
rect 6389 32027 6390 32325
rect 200 32026 6390 32027
rect 200 1000 500 32026
rect 9800 30570 10100 44430
rect 9800 30569 14534 30570
rect 9800 30271 14235 30569
rect 14533 30271 14534 30569
rect 9800 30270 14534 30271
rect 9800 1000 10100 30270
rect 24766 29497 29146 29498
rect 24766 29223 24767 29497
rect 25041 29223 29146 29497
rect 24766 29222 29146 29223
rect 15047 11920 15362 11921
rect 15047 11607 15048 11920
rect 15361 11607 15362 11920
rect 15047 4687 15362 11607
rect 23630 6735 27103 6736
rect 23630 6444 23631 6735
rect 23922 6444 27103 6735
rect 23630 6443 27103 6444
rect 21609 5608 21932 5609
rect 21609 5287 21610 5608
rect 21931 5287 21932 5608
rect 15047 4372 18282 4687
rect 17967 1699 18282 4372
rect 21609 4325 21932 5287
rect 21609 4002 22702 4325
rect 22379 1955 22702 4002
rect 26810 3448 27103 6443
rect 28870 3596 29146 29222
rect 28870 3518 30486 3596
rect 31312 3518 31432 3532
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 1699
rect 22480 0 22600 1955
rect 26896 0 27016 3448
rect 28870 3398 31432 3518
rect 28870 3320 30486 3398
rect 31312 0 31432 3398
use CurrentTrigger  CurrentTrigger_0
timestamp 1717084777
transform 0 1 16424 -1 0 27672
box -854 1682 19074 10100
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>

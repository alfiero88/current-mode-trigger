magic
tech sky130A
magscale 1 2
timestamp 1716907293
<< error_p >>
rect -415 381 -353 387
rect -287 381 -225 387
rect -159 381 -97 387
rect -31 381 31 387
rect 97 381 159 387
rect 225 381 287 387
rect 353 381 415 387
rect -415 347 -403 381
rect -287 347 -275 381
rect -159 347 -147 381
rect -31 347 -19 381
rect 97 347 109 381
rect 225 347 237 381
rect 353 347 365 381
rect -415 341 -353 347
rect -287 341 -225 347
rect -159 341 -97 347
rect -31 341 31 347
rect 97 341 159 347
rect 225 341 287 347
rect 353 341 415 347
rect -415 -347 -353 -341
rect -287 -347 -225 -341
rect -159 -347 -97 -341
rect -31 -347 31 -341
rect 97 -347 159 -341
rect 225 -347 287 -341
rect 353 -347 415 -341
rect -415 -381 -403 -347
rect -287 -381 -275 -347
rect -159 -381 -147 -347
rect -31 -381 -19 -347
rect 97 -381 109 -347
rect 225 -381 237 -347
rect 353 -381 365 -347
rect -415 -387 -353 -381
rect -287 -387 -225 -381
rect -159 -387 -97 -381
rect -31 -387 31 -381
rect 97 -387 159 -381
rect 225 -387 287 -381
rect 353 -387 415 -381
<< nwell >>
rect -615 -519 615 519
<< pmoslvt >>
rect -419 -300 -349 300
rect -291 -300 -221 300
rect -163 -300 -93 300
rect -35 -300 35 300
rect 93 -300 163 300
rect 221 -300 291 300
rect 349 -300 419 300
<< pdiff >>
rect -477 288 -419 300
rect -477 -288 -465 288
rect -431 -288 -419 288
rect -477 -300 -419 -288
rect -349 288 -291 300
rect -349 -288 -337 288
rect -303 -288 -291 288
rect -349 -300 -291 -288
rect -221 288 -163 300
rect -221 -288 -209 288
rect -175 -288 -163 288
rect -221 -300 -163 -288
rect -93 288 -35 300
rect -93 -288 -81 288
rect -47 -288 -35 288
rect -93 -300 -35 -288
rect 35 288 93 300
rect 35 -288 47 288
rect 81 -288 93 288
rect 35 -300 93 -288
rect 163 288 221 300
rect 163 -288 175 288
rect 209 -288 221 288
rect 163 -300 221 -288
rect 291 288 349 300
rect 291 -288 303 288
rect 337 -288 349 288
rect 291 -300 349 -288
rect 419 288 477 300
rect 419 -288 431 288
rect 465 -288 477 288
rect 419 -300 477 -288
<< pdiffc >>
rect -465 -288 -431 288
rect -337 -288 -303 288
rect -209 -288 -175 288
rect -81 -288 -47 288
rect 47 -288 81 288
rect 175 -288 209 288
rect 303 -288 337 288
rect 431 -288 465 288
<< nsubdiff >>
rect -579 449 -483 483
rect 483 449 579 483
rect -579 387 -545 449
rect 545 387 579 449
rect -579 -449 -545 -387
rect 545 -449 579 -387
rect -579 -483 -483 -449
rect 483 -483 579 -449
<< nsubdiffcont >>
rect -483 449 483 483
rect -579 -387 -545 387
rect 545 -387 579 387
rect -483 -483 483 -449
<< poly >>
rect -419 381 -349 397
rect -419 347 -403 381
rect -365 347 -349 381
rect -419 300 -349 347
rect -291 381 -221 397
rect -291 347 -275 381
rect -237 347 -221 381
rect -291 300 -221 347
rect -163 381 -93 397
rect -163 347 -147 381
rect -109 347 -93 381
rect -163 300 -93 347
rect -35 381 35 397
rect -35 347 -19 381
rect 19 347 35 381
rect -35 300 35 347
rect 93 381 163 397
rect 93 347 109 381
rect 147 347 163 381
rect 93 300 163 347
rect 221 381 291 397
rect 221 347 237 381
rect 275 347 291 381
rect 221 300 291 347
rect 349 381 419 397
rect 349 347 365 381
rect 403 347 419 381
rect 349 300 419 347
rect -419 -347 -349 -300
rect -419 -381 -403 -347
rect -365 -381 -349 -347
rect -419 -397 -349 -381
rect -291 -347 -221 -300
rect -291 -381 -275 -347
rect -237 -381 -221 -347
rect -291 -397 -221 -381
rect -163 -347 -93 -300
rect -163 -381 -147 -347
rect -109 -381 -93 -347
rect -163 -397 -93 -381
rect -35 -347 35 -300
rect -35 -381 -19 -347
rect 19 -381 35 -347
rect -35 -397 35 -381
rect 93 -347 163 -300
rect 93 -381 109 -347
rect 147 -381 163 -347
rect 93 -397 163 -381
rect 221 -347 291 -300
rect 221 -381 237 -347
rect 275 -381 291 -347
rect 221 -397 291 -381
rect 349 -347 419 -300
rect 349 -381 365 -347
rect 403 -381 419 -347
rect 349 -397 419 -381
<< polycont >>
rect -403 347 -365 381
rect -275 347 -237 381
rect -147 347 -109 381
rect -19 347 19 381
rect 109 347 147 381
rect 237 347 275 381
rect 365 347 403 381
rect -403 -381 -365 -347
rect -275 -381 -237 -347
rect -147 -381 -109 -347
rect -19 -381 19 -347
rect 109 -381 147 -347
rect 237 -381 275 -347
rect 365 -381 403 -347
<< locali >>
rect -579 449 -483 483
rect 483 449 579 483
rect -579 387 -545 449
rect 545 387 579 449
rect -419 347 -403 381
rect -365 347 -349 381
rect -291 347 -275 381
rect -237 347 -221 381
rect -163 347 -147 381
rect -109 347 -93 381
rect -35 347 -19 381
rect 19 347 35 381
rect 93 347 109 381
rect 147 347 163 381
rect 221 347 237 381
rect 275 347 291 381
rect 349 347 365 381
rect 403 347 419 381
rect -465 288 -431 304
rect -465 -304 -431 -288
rect -337 288 -303 304
rect -337 -304 -303 -288
rect -209 288 -175 304
rect -209 -304 -175 -288
rect -81 288 -47 304
rect -81 -304 -47 -288
rect 47 288 81 304
rect 47 -304 81 -288
rect 175 288 209 304
rect 175 -304 209 -288
rect 303 288 337 304
rect 303 -304 337 -288
rect 431 288 465 304
rect 431 -304 465 -288
rect -419 -381 -403 -347
rect -365 -381 -349 -347
rect -291 -381 -275 -347
rect -237 -381 -221 -347
rect -163 -381 -147 -347
rect -109 -381 -93 -347
rect -35 -381 -19 -347
rect 19 -381 35 -347
rect 93 -381 109 -347
rect 147 -381 163 -347
rect 221 -381 237 -347
rect 275 -381 291 -347
rect 349 -381 365 -347
rect 403 -381 419 -347
rect -579 -449 -545 -387
rect 545 -449 579 -387
rect -579 -483 -483 -449
rect 483 -483 579 -449
<< viali >>
rect -403 347 -365 381
rect -275 347 -237 381
rect -147 347 -109 381
rect -19 347 19 381
rect 109 347 147 381
rect 237 347 275 381
rect 365 347 403 381
rect -465 -288 -431 288
rect -337 -288 -303 288
rect -209 -288 -175 288
rect -81 -288 -47 288
rect 47 -288 81 288
rect 175 -288 209 288
rect 303 -288 337 288
rect 431 -288 465 288
rect -403 -381 -365 -347
rect -275 -381 -237 -347
rect -147 -381 -109 -347
rect -19 -381 19 -347
rect 109 -381 147 -347
rect 237 -381 275 -347
rect 365 -381 403 -347
<< metal1 >>
rect -415 381 -353 387
rect -415 347 -403 381
rect -365 347 -353 381
rect -415 341 -353 347
rect -287 381 -225 387
rect -287 347 -275 381
rect -237 347 -225 381
rect -287 341 -225 347
rect -159 381 -97 387
rect -159 347 -147 381
rect -109 347 -97 381
rect -159 341 -97 347
rect -31 381 31 387
rect -31 347 -19 381
rect 19 347 31 381
rect -31 341 31 347
rect 97 381 159 387
rect 97 347 109 381
rect 147 347 159 381
rect 97 341 159 347
rect 225 381 287 387
rect 225 347 237 381
rect 275 347 287 381
rect 225 341 287 347
rect 353 381 415 387
rect 353 347 365 381
rect 403 347 415 381
rect 353 341 415 347
rect -471 288 -425 300
rect -471 -288 -465 288
rect -431 -288 -425 288
rect -471 -300 -425 -288
rect -343 288 -297 300
rect -343 -288 -337 288
rect -303 -288 -297 288
rect -343 -300 -297 -288
rect -215 288 -169 300
rect -215 -288 -209 288
rect -175 -288 -169 288
rect -215 -300 -169 -288
rect -87 288 -41 300
rect -87 -288 -81 288
rect -47 -288 -41 288
rect -87 -300 -41 -288
rect 41 288 87 300
rect 41 -288 47 288
rect 81 -288 87 288
rect 41 -300 87 -288
rect 169 288 215 300
rect 169 -288 175 288
rect 209 -288 215 288
rect 169 -300 215 -288
rect 297 288 343 300
rect 297 -288 303 288
rect 337 -288 343 288
rect 297 -300 343 -288
rect 425 288 471 300
rect 425 -288 431 288
rect 465 -288 471 288
rect 425 -300 471 -288
rect -415 -347 -353 -341
rect -415 -381 -403 -347
rect -365 -381 -353 -347
rect -415 -387 -353 -381
rect -287 -347 -225 -341
rect -287 -381 -275 -347
rect -237 -381 -225 -347
rect -287 -387 -225 -381
rect -159 -347 -97 -341
rect -159 -381 -147 -347
rect -109 -381 -97 -347
rect -159 -387 -97 -381
rect -31 -347 31 -341
rect -31 -381 -19 -347
rect 19 -381 31 -347
rect -31 -387 31 -381
rect 97 -347 159 -341
rect 97 -381 109 -347
rect 147 -381 159 -347
rect 97 -387 159 -381
rect 225 -347 287 -341
rect 225 -381 237 -347
rect 275 -381 287 -347
rect 225 -387 287 -381
rect 353 -347 415 -341
rect 353 -381 365 -347
rect 403 -381 415 -347
rect 353 -387 415 -381
<< properties >>
string FIXED_BBOX -562 -466 562 466
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 3.0 l 0.35 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1717163641
<< metal1 >>
rect 28992 28608 29365 28645
rect 28992 28308 29028 28608
rect 29328 28308 29365 28608
rect 17380 26842 17680 26848
rect 21380 26845 21736 26870
rect 20593 26842 21736 26845
rect 17680 26542 21736 26842
rect 17380 26536 17680 26542
rect 20593 26539 21736 26542
rect 21380 24456 21736 26539
rect 25472 25938 27587 26005
rect 25472 25818 27400 25938
rect 27520 25818 27587 25938
rect 25472 25752 27587 25818
rect 25472 24566 25725 25752
rect 28992 24362 29365 28308
rect 22324 12894 23474 12967
rect 22324 12774 22396 12894
rect 22516 12774 23474 12894
rect 22324 12702 23474 12774
rect 26769 6076 27003 6879
rect 26769 5956 26826 6076
rect 26946 5956 27003 6076
rect 26769 5899 27003 5956
rect 24775 4064 25009 5425
rect 24775 3944 24832 4064
rect 24952 3944 25009 4064
rect 24775 3887 25009 3944
<< via1 >>
rect 29028 28308 29328 28608
rect 17380 26542 17680 26842
rect 27400 25818 27520 25938
rect 22396 12774 22516 12894
rect 26826 5956 26946 6076
rect 24832 3944 24952 4064
<< metal2 >>
rect 19297 28608 19587 28612
rect 19292 28603 29028 28608
rect 19292 28313 19297 28603
rect 19587 28313 29028 28603
rect 19292 28308 29028 28313
rect 29328 28308 29334 28608
rect 19297 28304 19587 28308
rect 15387 26842 15677 26846
rect 15382 26837 17380 26842
rect 15382 26547 15387 26837
rect 15677 26547 17380 26837
rect 15382 26542 17380 26547
rect 17680 26542 17686 26842
rect 15387 26538 15677 26542
rect 27394 25818 27400 25938
rect 27520 25818 31432 25938
rect 31312 20597 31432 25818
rect 31308 20487 31317 20597
rect 31427 20487 31436 20597
rect 31312 20482 31432 20487
rect 18064 12774 22396 12894
rect 22516 12774 22522 12894
rect 18064 7481 18184 12774
rect 18060 7371 18069 7481
rect 18179 7371 18188 7481
rect 18064 7366 18184 7371
rect 26826 6076 26946 6082
rect 26826 5786 26946 5956
rect 26826 5666 27016 5786
rect 24832 4064 24952 4070
rect 24832 2581 24952 3944
rect 26896 3191 27016 5666
rect 26892 3081 26901 3191
rect 27011 3081 27020 3191
rect 26896 3076 27016 3081
rect 24828 2471 24837 2581
rect 24947 2471 24956 2581
rect 24832 2466 24952 2471
<< via2 >>
rect 19297 28313 19587 28603
rect 15387 26547 15677 26837
rect 31317 20487 31427 20597
rect 18069 7371 18179 7481
rect 26901 3081 27011 3191
rect 24837 2471 24947 2581
<< metal3 >>
rect 5937 28608 6235 28613
rect 5936 28607 19592 28608
rect 5936 28309 5937 28607
rect 6235 28603 19592 28607
rect 6235 28313 19297 28603
rect 19587 28313 19592 28603
rect 6235 28309 19592 28313
rect 5936 28308 19592 28309
rect 5937 28303 6235 28308
rect 13963 26842 14261 26847
rect 13962 26841 15682 26842
rect 13962 26543 13963 26841
rect 14261 26837 15682 26841
rect 14261 26547 15387 26837
rect 15677 26547 15682 26837
rect 14261 26543 15682 26547
rect 13962 26542 15682 26543
rect 13963 26537 14261 26542
rect 31312 20597 31432 20602
rect 31312 20487 31317 20597
rect 31427 20487 31432 20597
rect 31312 9489 31432 20487
rect 31307 9371 31313 9489
rect 31431 9371 31437 9489
rect 31312 9370 31432 9371
rect 18064 7481 18184 7486
rect 18064 7371 18069 7481
rect 18179 7371 18184 7481
rect 18064 4583 18184 7371
rect 18059 4465 18065 4583
rect 18183 4465 18189 4583
rect 18064 4464 18184 4465
rect 26896 3191 27016 3196
rect 26896 3081 26901 3191
rect 27011 3081 27016 3191
rect 24832 2581 24952 2586
rect 24832 2471 24837 2581
rect 24947 2471 24952 2581
rect 23557 2210 23675 2215
rect 24832 2210 24952 2471
rect 26896 2253 27016 3081
rect 23556 2209 24952 2210
rect 23556 2091 23557 2209
rect 23675 2091 24952 2209
rect 26891 2135 26897 2253
rect 27015 2135 27021 2253
rect 26896 2134 27016 2135
rect 23556 2090 24952 2091
rect 23557 2085 23675 2090
<< via3 >>
rect 5937 28309 6235 28607
rect 13963 26543 14261 26841
rect 31313 9371 31431 9489
rect 18065 4465 18183 4583
rect 23557 2091 23675 2209
rect 26897 2135 27015 2253
<< metal4 >>
rect 798 44838 858 45152
rect 1534 44838 1594 45152
rect 2270 44838 2330 45152
rect 3006 44838 3066 45152
rect 3742 44838 3802 45152
rect 4478 44838 4538 45152
rect 5214 44838 5274 45152
rect 5950 44838 6010 45152
rect 6686 44838 6746 45152
rect 7422 44838 7482 45152
rect 8158 44838 8218 45152
rect 8894 44838 8954 45152
rect 9630 44838 9690 45152
rect 10366 44838 10426 45152
rect 11102 44838 11162 45152
rect 11838 44838 11898 45152
rect 12574 44838 12634 45152
rect 13310 44838 13370 45152
rect 14046 44838 14106 45152
rect 14782 44838 14842 45152
rect 15518 44838 15578 45152
rect 16254 44838 16314 45152
rect 16990 44838 17050 45152
rect 17726 44838 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 632 44488 17862 44838
rect 200 28608 500 44152
rect 200 28607 6236 28608
rect 200 28309 5937 28607
rect 6235 28309 6236 28607
rect 200 28308 6236 28309
rect 200 1000 500 28308
rect 9800 26842 10100 44488
rect 9800 26841 14262 26842
rect 9800 26543 13963 26841
rect 14261 26543 14262 26841
rect 9800 26542 14262 26543
rect 9800 1000 10100 26542
rect 31312 9489 31432 9490
rect 31312 9371 31313 9489
rect 31431 9371 31432 9489
rect 18064 4583 18184 4584
rect 18064 4465 18065 4583
rect 18183 4465 18184 4583
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 4465
rect 26896 2253 27016 2254
rect 22480 2209 23676 2210
rect 22480 2091 23557 2209
rect 23675 2091 23676 2209
rect 22480 2090 23676 2091
rect 26896 2135 26897 2253
rect 27015 2135 27016 2253
rect 22480 0 22600 2090
rect 26896 0 27016 2135
rect 31312 0 31432 9371
use CurrentTrigger  CurrentTrigger_0
timestamp 1717084777
transform 0 1 19520 -1 0 24076
box -854 1682 19074 10100
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 4800 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 4800 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1716907293
<< error_p >>
rect -159 248 -97 254
rect -31 248 31 254
rect 97 248 159 254
rect -159 214 -147 248
rect -31 214 -19 248
rect 97 214 109 248
rect -159 208 -97 214
rect -31 208 31 214
rect 97 208 159 214
rect -159 -214 -97 -208
rect -31 -214 31 -208
rect 97 -214 159 -208
rect -159 -248 -147 -214
rect -31 -248 -19 -214
rect 97 -248 109 -214
rect -159 -254 -97 -248
rect -31 -254 31 -248
rect 97 -254 159 -248
<< nwell >>
rect -359 -386 359 386
<< pmoslvt >>
rect -163 -167 -93 167
rect -35 -167 35 167
rect 93 -167 163 167
<< pdiff >>
rect -221 155 -163 167
rect -221 -155 -209 155
rect -175 -155 -163 155
rect -221 -167 -163 -155
rect -93 155 -35 167
rect -93 -155 -81 155
rect -47 -155 -35 155
rect -93 -167 -35 -155
rect 35 155 93 167
rect 35 -155 47 155
rect 81 -155 93 155
rect 35 -167 93 -155
rect 163 155 221 167
rect 163 -155 175 155
rect 209 -155 221 155
rect 163 -167 221 -155
<< pdiffc >>
rect -209 -155 -175 155
rect -81 -155 -47 155
rect 47 -155 81 155
rect 175 -155 209 155
<< nsubdiff >>
rect -323 316 -227 350
rect 227 316 323 350
rect -323 254 -289 316
rect 289 254 323 316
rect -323 -316 -289 -254
rect 289 -316 323 -254
rect -323 -350 -227 -316
rect 227 -350 323 -316
<< nsubdiffcont >>
rect -227 316 227 350
rect -323 -254 -289 254
rect 289 -254 323 254
rect -227 -350 227 -316
<< poly >>
rect -163 248 -93 264
rect -163 214 -147 248
rect -109 214 -93 248
rect -163 167 -93 214
rect -35 248 35 264
rect -35 214 -19 248
rect 19 214 35 248
rect -35 167 35 214
rect 93 248 163 264
rect 93 214 109 248
rect 147 214 163 248
rect 93 167 163 214
rect -163 -214 -93 -167
rect -163 -248 -147 -214
rect -109 -248 -93 -214
rect -163 -264 -93 -248
rect -35 -214 35 -167
rect -35 -248 -19 -214
rect 19 -248 35 -214
rect -35 -264 35 -248
rect 93 -214 163 -167
rect 93 -248 109 -214
rect 147 -248 163 -214
rect 93 -264 163 -248
<< polycont >>
rect -147 214 -109 248
rect -19 214 19 248
rect 109 214 147 248
rect -147 -248 -109 -214
rect -19 -248 19 -214
rect 109 -248 147 -214
<< locali >>
rect -323 316 -227 350
rect 227 316 323 350
rect -323 254 -289 316
rect 289 254 323 316
rect -163 214 -147 248
rect -109 214 -93 248
rect -35 214 -19 248
rect 19 214 35 248
rect 93 214 109 248
rect 147 214 163 248
rect -209 155 -175 171
rect -209 -171 -175 -155
rect -81 155 -47 171
rect -81 -171 -47 -155
rect 47 155 81 171
rect 47 -171 81 -155
rect 175 155 209 171
rect 175 -171 209 -155
rect -163 -248 -147 -214
rect -109 -248 -93 -214
rect -35 -248 -19 -214
rect 19 -248 35 -214
rect 93 -248 109 -214
rect 147 -248 163 -214
rect -323 -316 -289 -254
rect 289 -316 323 -254
rect -323 -350 -227 -316
rect 227 -350 323 -316
<< viali >>
rect -147 214 -109 248
rect -19 214 19 248
rect 109 214 147 248
rect -209 -155 -175 155
rect -81 -155 -47 155
rect 47 -155 81 155
rect 175 -155 209 155
rect -147 -248 -109 -214
rect -19 -248 19 -214
rect 109 -248 147 -214
<< metal1 >>
rect -159 248 -97 254
rect -159 214 -147 248
rect -109 214 -97 248
rect -159 208 -97 214
rect -31 248 31 254
rect -31 214 -19 248
rect 19 214 31 248
rect -31 208 31 214
rect 97 248 159 254
rect 97 214 109 248
rect 147 214 159 248
rect 97 208 159 214
rect -215 155 -169 167
rect -215 -155 -209 155
rect -175 -155 -169 155
rect -215 -167 -169 -155
rect -87 155 -41 167
rect -87 -155 -81 155
rect -47 -155 -41 155
rect -87 -167 -41 -155
rect 41 155 87 167
rect 41 -155 47 155
rect 81 -155 87 155
rect 41 -167 87 -155
rect 169 155 215 167
rect 169 -155 175 155
rect 209 -155 215 155
rect 169 -167 215 -155
rect -159 -214 -97 -208
rect -159 -248 -147 -214
rect -109 -248 -97 -214
rect -159 -254 -97 -248
rect -31 -214 31 -208
rect -31 -248 -19 -214
rect 19 -248 31 -214
rect -31 -254 31 -248
rect 97 -214 159 -208
rect 97 -248 109 -214
rect 147 -248 159 -214
rect 97 -254 159 -248
<< properties >>
string FIXED_BBOX -306 -333 306 333
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1.6666666666666667 l 0.35 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

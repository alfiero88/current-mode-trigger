magic
tech sky130A
timestamp 1716907293
<< pwell >>
rect -427 -155 427 155
<< nmoslvt >>
rect -329 -50 -129 50
rect -100 -50 100 50
rect 129 -50 329 50
<< ndiff >>
rect -358 44 -329 50
rect -358 -44 -352 44
rect -335 -44 -329 44
rect -358 -50 -329 -44
rect -129 44 -100 50
rect -129 -44 -123 44
rect -106 -44 -100 44
rect -129 -50 -100 -44
rect 100 44 129 50
rect 100 -44 106 44
rect 123 -44 129 44
rect 100 -50 129 -44
rect 329 44 358 50
rect 329 -44 335 44
rect 352 -44 358 44
rect 329 -50 358 -44
<< ndiffc >>
rect -352 -44 -335 44
rect -123 -44 -106 44
rect 106 -44 123 44
rect 335 -44 352 44
<< psubdiff >>
rect -409 120 -361 137
rect 361 120 409 137
rect -409 89 -392 120
rect 392 89 409 120
rect -409 -120 -392 -89
rect 392 -120 409 -89
rect -409 -137 -361 -120
rect 361 -137 409 -120
<< psubdiffcont >>
rect -361 120 361 137
rect -409 -89 -392 89
rect 392 -89 409 89
rect -361 -137 361 -120
<< poly >>
rect -329 86 -129 94
rect -329 69 -321 86
rect -137 69 -129 86
rect -329 50 -129 69
rect -100 86 100 94
rect -100 69 -92 86
rect 92 69 100 86
rect -100 50 100 69
rect 129 86 329 94
rect 129 69 137 86
rect 321 69 329 86
rect 129 50 329 69
rect -329 -69 -129 -50
rect -329 -86 -321 -69
rect -137 -86 -129 -69
rect -329 -94 -129 -86
rect -100 -69 100 -50
rect -100 -86 -92 -69
rect 92 -86 100 -69
rect -100 -94 100 -86
rect 129 -69 329 -50
rect 129 -86 137 -69
rect 321 -86 329 -69
rect 129 -94 329 -86
<< polycont >>
rect -321 69 -137 86
rect -92 69 92 86
rect 137 69 321 86
rect -321 -86 -137 -69
rect -92 -86 92 -69
rect 137 -86 321 -69
<< locali >>
rect -409 120 -361 137
rect 361 120 409 137
rect -409 89 -392 120
rect 392 89 409 120
rect -329 69 -321 86
rect -137 69 -129 86
rect -100 69 -92 86
rect 92 69 100 86
rect 129 69 137 86
rect 321 69 329 86
rect -352 44 -335 52
rect -352 -52 -335 -44
rect -123 44 -106 52
rect -123 -52 -106 -44
rect 106 44 123 52
rect 106 -52 123 -44
rect 335 44 352 52
rect 335 -52 352 -44
rect -329 -86 -321 -69
rect -137 -86 -129 -69
rect -100 -86 -92 -69
rect 92 -86 100 -69
rect 129 -86 137 -69
rect 321 -86 329 -69
rect -409 -120 -392 -89
rect 392 -120 409 -89
rect -409 -137 -361 -120
rect 361 -137 409 -120
<< viali >>
rect -321 69 -137 86
rect -92 69 92 86
rect 137 69 321 86
rect -352 -44 -335 44
rect -123 -44 -106 44
rect 106 -44 123 44
rect 335 -44 352 44
rect -321 -86 -137 -69
rect -92 -86 92 -69
rect 137 -86 321 -69
<< metal1 >>
rect -327 86 -131 89
rect -327 69 -321 86
rect -137 69 -131 86
rect -327 66 -131 69
rect -98 86 98 89
rect -98 69 -92 86
rect 92 69 98 86
rect -98 66 98 69
rect 131 86 327 89
rect 131 69 137 86
rect 321 69 327 86
rect 131 66 327 69
rect -355 44 -332 50
rect -355 -44 -352 44
rect -335 -44 -332 44
rect -355 -50 -332 -44
rect -126 44 -103 50
rect -126 -44 -123 44
rect -106 -44 -103 44
rect -126 -50 -103 -44
rect 103 44 126 50
rect 103 -44 106 44
rect 123 -44 126 44
rect 103 -50 126 -44
rect 332 44 355 50
rect 332 -44 335 44
rect 352 -44 355 44
rect 332 -50 355 -44
rect -327 -69 -131 -66
rect -327 -86 -321 -69
rect -137 -86 -131 -69
rect -327 -89 -131 -86
rect -98 -69 98 -66
rect -98 -86 -92 -69
rect 92 -86 98 -69
rect -98 -89 98 -86
rect 131 -69 327 -66
rect 131 -86 137 -69
rect 321 -86 327 -69
rect 131 -89 327 -86
<< properties >>
string FIXED_BBOX -400 -128 400 128
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.0 l 2.0 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

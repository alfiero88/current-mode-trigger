VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_alfiero88_CurrentTrigger
  CLASS BLOCK ;
  FOREIGN tt_um_alfiero88_CurrentTrigger ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.350000 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.000000 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.530000 ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 10.312400 ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 95.610 132.920 100.710 137.880 ;
        RECT 105.270 132.850 110.370 137.880 ;
      LAYER nwell ;
        RECT 114.400 131.730 119.590 137.880 ;
        RECT 122.790 132.810 127.980 137.770 ;
      LAYER pwell ;
        RECT 96.190 111.170 102.290 122.710 ;
        RECT 96.250 95.570 102.350 107.110 ;
      LAYER nwell ;
        RECT 107.020 99.570 110.710 119.060 ;
        RECT 114.850 99.570 118.540 119.060 ;
      LAYER pwell ;
        RECT 99.240 86.420 102.340 91.960 ;
      LAYER nwell ;
        RECT 112.380 86.320 116.710 92.470 ;
        RECT 122.690 84.410 126.880 115.690 ;
      LAYER pwell ;
        RECT 99.270 72.450 102.370 77.990 ;
        RECT 113.510 70.900 116.610 79.440 ;
      LAYER nwell ;
        RECT 122.340 75.020 126.200 78.610 ;
      LAYER pwell ;
        RECT 105.040 62.460 108.140 64.570 ;
      LAYER nwell ;
        RECT 110.370 62.310 114.560 64.620 ;
      LAYER pwell ;
        RECT 105.040 57.260 108.640 59.890 ;
      LAYER nwell ;
        RECT 110.370 56.890 114.560 60.480 ;
      LAYER pwell ;
        RECT 103.600 49.950 108.700 53.060 ;
      LAYER nwell ;
        RECT 110.370 48.750 115.560 54.260 ;
        RECT 122.140 48.640 126.330 70.050 ;
      LAYER li1 ;
        RECT 105.900 137.700 109.750 137.750 ;
        RECT 115.040 137.700 118.940 137.730 ;
        RECT 95.790 137.530 100.530 137.700 ;
        RECT 95.790 137.250 95.960 137.530 ;
        RECT 95.750 133.560 95.960 137.250 ;
        RECT 96.640 136.960 99.680 137.130 ;
        RECT 96.300 133.900 96.470 136.900 ;
        RECT 99.850 133.900 100.020 136.900 ;
        RECT 96.640 133.670 99.680 133.840 ;
        RECT 95.790 133.270 95.960 133.560 ;
        RECT 100.360 133.270 100.530 137.530 ;
        RECT 95.790 133.100 100.530 133.270 ;
        RECT 105.450 137.530 110.190 137.700 ;
        RECT 105.450 133.200 105.620 137.530 ;
        RECT 105.960 136.640 106.130 136.970 ;
        RECT 106.300 136.960 109.340 137.130 ;
        RECT 106.300 136.480 109.340 136.650 ;
        RECT 105.960 135.680 106.130 136.010 ;
        RECT 106.300 136.000 109.340 136.170 ;
        RECT 109.510 136.160 109.680 136.490 ;
        RECT 106.300 135.520 109.340 135.690 ;
        RECT 105.960 134.720 106.130 135.050 ;
        RECT 106.300 135.040 109.340 135.210 ;
        RECT 109.510 135.200 109.680 135.530 ;
        RECT 106.300 134.560 109.340 134.730 ;
        RECT 105.960 133.760 106.130 134.090 ;
        RECT 106.300 134.080 109.340 134.250 ;
        RECT 109.510 134.240 109.680 134.570 ;
        RECT 106.300 133.600 109.340 133.770 ;
        RECT 110.020 133.200 110.190 137.530 ;
        RECT 105.450 133.030 110.190 133.200 ;
        RECT 114.580 137.530 119.410 137.700 ;
        RECT 114.580 132.080 114.750 137.530 ;
        RECT 115.475 136.960 118.515 137.130 ;
        RECT 115.090 136.550 115.260 136.900 ;
        RECT 118.730 136.550 118.900 136.900 ;
        RECT 115.475 136.320 118.515 136.490 ;
        RECT 115.090 135.910 115.260 136.260 ;
        RECT 118.730 135.910 118.900 136.260 ;
        RECT 115.475 135.680 118.515 135.850 ;
        RECT 115.090 135.270 115.260 135.620 ;
        RECT 118.730 135.270 118.900 135.620 ;
        RECT 115.475 135.040 118.515 135.210 ;
        RECT 115.090 134.630 115.260 134.980 ;
        RECT 118.730 134.630 118.900 134.980 ;
        RECT 115.475 134.400 118.515 134.570 ;
        RECT 115.090 133.990 115.260 134.340 ;
        RECT 118.730 133.990 118.900 134.340 ;
        RECT 115.475 133.760 118.515 133.930 ;
        RECT 115.090 133.350 115.260 133.700 ;
        RECT 118.730 133.350 118.900 133.700 ;
        RECT 115.475 133.120 118.515 133.290 ;
        RECT 115.090 132.710 115.260 133.060 ;
        RECT 118.730 132.710 118.900 133.060 ;
        RECT 115.475 132.480 118.515 132.650 ;
        RECT 119.240 132.080 119.410 137.530 ;
        RECT 122.970 137.420 127.800 137.590 ;
        RECT 122.970 133.160 123.140 137.420 ;
        RECT 127.630 137.130 127.800 137.420 ;
        RECT 123.865 136.850 126.905 137.020 ;
        RECT 123.480 133.790 123.650 136.790 ;
        RECT 127.120 133.790 127.290 136.790 ;
        RECT 123.865 133.560 126.905 133.730 ;
        RECT 127.630 133.450 127.830 137.130 ;
        RECT 127.630 133.160 127.800 133.450 ;
        RECT 122.970 132.990 127.800 133.160 ;
        RECT 114.580 131.910 119.410 132.080 ;
        RECT 96.370 122.360 102.110 122.530 ;
        RECT 96.370 122.080 96.540 122.360 ;
        RECT 96.300 111.800 96.540 122.080 ;
        RECT 97.220 121.790 101.260 121.960 ;
        RECT 96.880 118.730 97.050 121.730 ;
        RECT 101.430 118.730 101.600 121.730 ;
        RECT 97.220 118.500 101.260 118.670 ;
        RECT 96.880 115.440 97.050 118.440 ;
        RECT 101.430 115.440 101.600 118.440 ;
        RECT 97.220 115.210 101.260 115.380 ;
        RECT 96.880 112.150 97.050 115.150 ;
        RECT 101.430 112.150 101.600 115.150 ;
        RECT 97.220 111.920 101.260 112.090 ;
        RECT 96.370 111.520 96.540 111.800 ;
        RECT 101.940 111.520 102.110 122.360 ;
        RECT 96.370 111.350 102.110 111.520 ;
        RECT 107.200 118.710 110.530 118.880 ;
        RECT 96.430 106.760 102.170 106.930 ;
        RECT 96.430 106.470 96.600 106.760 ;
        RECT 96.360 96.210 96.600 106.470 ;
        RECT 97.280 106.190 101.320 106.360 ;
        RECT 96.940 103.130 97.110 106.130 ;
        RECT 101.490 103.130 101.660 106.130 ;
        RECT 97.280 102.900 101.320 103.070 ;
        RECT 96.940 99.840 97.110 102.840 ;
        RECT 101.490 99.840 101.660 102.840 ;
        RECT 97.280 99.610 101.320 99.780 ;
        RECT 96.940 96.550 97.110 99.550 ;
        RECT 101.490 96.550 101.660 99.550 ;
        RECT 97.280 96.320 101.320 96.490 ;
        RECT 96.430 95.920 96.600 96.210 ;
        RECT 102.000 95.920 102.170 106.760 ;
        RECT 107.200 99.920 107.370 118.710 ;
        RECT 110.360 118.450 110.530 118.710 ;
        RECT 115.030 118.710 118.360 118.880 ;
        RECT 108.095 118.140 109.635 118.310 ;
        RECT 107.710 117.380 107.880 118.080 ;
        RECT 109.850 117.380 110.020 118.080 ;
        RECT 108.095 117.150 109.635 117.320 ;
        RECT 107.710 116.390 107.880 117.090 ;
        RECT 109.850 116.390 110.020 117.090 ;
        RECT 108.095 116.160 109.635 116.330 ;
        RECT 107.710 115.400 107.880 116.100 ;
        RECT 109.850 115.400 110.020 116.100 ;
        RECT 108.095 115.170 109.635 115.340 ;
        RECT 107.710 114.410 107.880 115.110 ;
        RECT 109.850 114.410 110.020 115.110 ;
        RECT 108.095 114.180 109.635 114.350 ;
        RECT 107.710 113.420 107.880 114.120 ;
        RECT 109.850 113.420 110.020 114.120 ;
        RECT 108.095 113.190 109.635 113.360 ;
        RECT 107.710 112.430 107.880 113.130 ;
        RECT 109.850 112.430 110.020 113.130 ;
        RECT 108.095 112.200 109.635 112.370 ;
        RECT 107.710 111.440 107.880 112.140 ;
        RECT 109.850 111.440 110.020 112.140 ;
        RECT 108.095 111.210 109.635 111.380 ;
        RECT 107.710 110.450 107.880 111.150 ;
        RECT 109.850 110.450 110.020 111.150 ;
        RECT 108.095 110.220 109.635 110.390 ;
        RECT 107.710 109.460 107.880 110.160 ;
        RECT 109.850 109.460 110.020 110.160 ;
        RECT 108.095 109.230 109.635 109.400 ;
        RECT 107.710 108.470 107.880 109.170 ;
        RECT 109.850 108.470 110.020 109.170 ;
        RECT 108.095 108.240 109.635 108.410 ;
        RECT 107.710 107.480 107.880 108.180 ;
        RECT 109.850 107.480 110.020 108.180 ;
        RECT 108.095 107.250 109.635 107.420 ;
        RECT 107.710 106.490 107.880 107.190 ;
        RECT 109.850 106.490 110.020 107.190 ;
        RECT 108.095 106.260 109.635 106.430 ;
        RECT 107.710 105.500 107.880 106.200 ;
        RECT 109.850 105.500 110.020 106.200 ;
        RECT 108.095 105.270 109.635 105.440 ;
        RECT 107.710 104.510 107.880 105.210 ;
        RECT 109.850 104.510 110.020 105.210 ;
        RECT 108.095 104.280 109.635 104.450 ;
        RECT 107.710 103.520 107.880 104.220 ;
        RECT 109.850 103.520 110.020 104.220 ;
        RECT 108.095 103.290 109.635 103.460 ;
        RECT 107.710 102.530 107.880 103.230 ;
        RECT 109.850 102.530 110.020 103.230 ;
        RECT 108.095 102.300 109.635 102.470 ;
        RECT 107.710 101.540 107.880 102.240 ;
        RECT 109.850 101.540 110.020 102.240 ;
        RECT 108.095 101.310 109.635 101.480 ;
        RECT 107.710 100.550 107.880 101.250 ;
        RECT 109.850 100.550 110.020 101.250 ;
        RECT 108.095 100.320 109.635 100.490 ;
        RECT 110.360 100.180 110.770 118.450 ;
        RECT 110.360 99.920 110.530 100.180 ;
        RECT 107.200 99.750 110.530 99.920 ;
        RECT 115.030 99.920 115.200 118.710 ;
        RECT 118.190 118.310 118.360 118.710 ;
        RECT 115.925 118.140 117.465 118.310 ;
        RECT 115.540 117.380 115.710 118.080 ;
        RECT 117.680 117.380 117.850 118.080 ;
        RECT 115.925 117.150 117.465 117.320 ;
        RECT 115.540 116.390 115.710 117.090 ;
        RECT 117.680 116.390 117.850 117.090 ;
        RECT 115.925 116.160 117.465 116.330 ;
        RECT 115.540 115.400 115.710 116.100 ;
        RECT 117.680 115.400 117.850 116.100 ;
        RECT 115.925 115.170 117.465 115.340 ;
        RECT 115.540 114.410 115.710 115.110 ;
        RECT 117.680 114.410 117.850 115.110 ;
        RECT 115.925 114.180 117.465 114.350 ;
        RECT 115.540 113.420 115.710 114.120 ;
        RECT 117.680 113.420 117.850 114.120 ;
        RECT 115.925 113.190 117.465 113.360 ;
        RECT 115.540 112.430 115.710 113.130 ;
        RECT 117.680 112.430 117.850 113.130 ;
        RECT 115.925 112.200 117.465 112.370 ;
        RECT 115.540 111.440 115.710 112.140 ;
        RECT 117.680 111.440 117.850 112.140 ;
        RECT 115.925 111.210 117.465 111.380 ;
        RECT 115.540 110.450 115.710 111.150 ;
        RECT 117.680 110.450 117.850 111.150 ;
        RECT 115.925 110.220 117.465 110.390 ;
        RECT 115.540 109.460 115.710 110.160 ;
        RECT 117.680 109.460 117.850 110.160 ;
        RECT 115.925 109.230 117.465 109.400 ;
        RECT 115.540 108.470 115.710 109.170 ;
        RECT 117.680 108.470 117.850 109.170 ;
        RECT 115.925 108.240 117.465 108.410 ;
        RECT 115.540 107.480 115.710 108.180 ;
        RECT 117.680 107.480 117.850 108.180 ;
        RECT 115.925 107.250 117.465 107.420 ;
        RECT 115.540 106.490 115.710 107.190 ;
        RECT 117.680 106.490 117.850 107.190 ;
        RECT 115.925 106.260 117.465 106.430 ;
        RECT 115.540 105.500 115.710 106.200 ;
        RECT 117.680 105.500 117.850 106.200 ;
        RECT 115.925 105.270 117.465 105.440 ;
        RECT 115.540 104.510 115.710 105.210 ;
        RECT 117.680 104.510 117.850 105.210 ;
        RECT 115.925 104.280 117.465 104.450 ;
        RECT 115.540 103.520 115.710 104.220 ;
        RECT 117.680 103.520 117.850 104.220 ;
        RECT 115.925 103.290 117.465 103.460 ;
        RECT 115.540 102.530 115.710 103.230 ;
        RECT 117.680 102.530 117.850 103.230 ;
        RECT 115.925 102.300 117.465 102.470 ;
        RECT 115.540 101.540 115.710 102.240 ;
        RECT 117.680 101.540 117.850 102.240 ;
        RECT 115.925 101.310 117.465 101.480 ;
        RECT 115.540 100.550 115.710 101.250 ;
        RECT 117.680 100.550 117.850 101.250 ;
        RECT 115.925 100.320 117.465 100.490 ;
        RECT 118.180 100.210 118.480 118.310 ;
        RECT 122.870 115.340 126.700 115.510 ;
        RECT 118.190 99.920 118.360 100.210 ;
        RECT 115.030 99.750 118.360 99.920 ;
        RECT 96.430 95.750 102.170 95.920 ;
        RECT 112.560 92.120 116.530 92.290 ;
        RECT 99.420 91.610 102.160 91.780 ;
        RECT 99.420 91.340 99.590 91.610 ;
        RECT 99.360 87.040 99.590 91.340 ;
        RECT 100.270 91.040 101.310 91.210 ;
        RECT 99.930 89.980 100.100 90.980 ;
        RECT 101.480 89.980 101.650 90.980 ;
        RECT 100.270 89.750 101.310 89.920 ;
        RECT 99.930 88.690 100.100 89.690 ;
        RECT 101.480 88.690 101.650 89.690 ;
        RECT 100.270 88.460 101.310 88.630 ;
        RECT 99.930 87.400 100.100 88.400 ;
        RECT 101.480 87.400 101.650 88.400 ;
        RECT 100.270 87.170 101.310 87.340 ;
        RECT 99.420 86.770 99.590 87.040 ;
        RECT 101.990 86.770 102.160 91.610 ;
        RECT 99.420 86.600 102.160 86.770 ;
        RECT 112.560 86.670 112.730 92.120 ;
        RECT 116.360 91.870 116.530 92.120 ;
        RECT 113.455 91.550 115.635 91.720 ;
        RECT 113.070 91.140 113.240 91.490 ;
        RECT 115.850 91.140 116.020 91.490 ;
        RECT 113.455 90.910 115.635 91.080 ;
        RECT 113.070 90.500 113.240 90.850 ;
        RECT 115.850 90.500 116.020 90.850 ;
        RECT 113.455 90.270 115.635 90.440 ;
        RECT 113.070 89.860 113.240 90.210 ;
        RECT 115.850 89.860 116.020 90.210 ;
        RECT 113.455 89.630 115.635 89.800 ;
        RECT 113.070 89.220 113.240 89.570 ;
        RECT 115.850 89.220 116.020 89.570 ;
        RECT 113.455 88.990 115.635 89.160 ;
        RECT 113.070 88.580 113.240 88.930 ;
        RECT 115.850 88.580 116.020 88.930 ;
        RECT 113.455 88.350 115.635 88.520 ;
        RECT 113.070 87.940 113.240 88.290 ;
        RECT 115.850 87.940 116.020 88.290 ;
        RECT 113.455 87.710 115.635 87.880 ;
        RECT 113.070 87.300 113.240 87.650 ;
        RECT 115.850 87.300 116.020 87.650 ;
        RECT 113.455 87.070 115.635 87.240 ;
        RECT 116.360 86.920 116.620 91.870 ;
        RECT 116.360 86.670 116.530 86.920 ;
        RECT 112.560 86.500 116.530 86.670 ;
        RECT 122.870 84.760 123.040 115.340 ;
        RECT 126.530 115.060 126.700 115.340 ;
        RECT 123.765 114.770 125.805 114.940 ;
        RECT 123.380 111.710 123.550 114.710 ;
        RECT 126.020 111.710 126.190 114.710 ;
        RECT 123.765 111.480 125.805 111.650 ;
        RECT 123.380 108.420 123.550 111.420 ;
        RECT 126.020 108.420 126.190 111.420 ;
        RECT 123.765 108.190 125.805 108.360 ;
        RECT 123.380 105.130 123.550 108.130 ;
        RECT 126.020 105.130 126.190 108.130 ;
        RECT 123.765 104.900 125.805 105.070 ;
        RECT 123.380 101.840 123.550 104.840 ;
        RECT 126.020 101.840 126.190 104.840 ;
        RECT 123.765 101.610 125.805 101.780 ;
        RECT 123.380 98.550 123.550 101.550 ;
        RECT 126.020 98.550 126.190 101.550 ;
        RECT 123.765 98.320 125.805 98.490 ;
        RECT 123.380 95.260 123.550 98.260 ;
        RECT 126.020 95.260 126.190 98.260 ;
        RECT 123.765 95.030 125.805 95.200 ;
        RECT 123.380 91.970 123.550 94.970 ;
        RECT 126.020 91.970 126.190 94.970 ;
        RECT 123.765 91.740 125.805 91.910 ;
        RECT 123.380 88.680 123.550 91.680 ;
        RECT 126.020 88.680 126.190 91.680 ;
        RECT 123.765 88.450 125.805 88.620 ;
        RECT 123.380 85.390 123.550 88.390 ;
        RECT 126.020 85.390 126.190 88.390 ;
        RECT 123.765 85.160 125.805 85.330 ;
        RECT 126.530 85.020 126.770 115.060 ;
        RECT 126.530 84.760 126.700 85.020 ;
        RECT 122.870 84.590 126.700 84.760 ;
        RECT 113.690 79.090 116.430 79.260 ;
        RECT 113.690 78.840 113.860 79.090 ;
        RECT 99.450 77.640 102.190 77.810 ;
        RECT 99.450 77.390 99.620 77.640 ;
        RECT 99.300 73.050 99.620 77.390 ;
        RECT 100.300 77.070 101.340 77.240 ;
        RECT 99.960 76.010 100.130 77.010 ;
        RECT 101.510 76.010 101.680 77.010 ;
        RECT 100.300 75.780 101.340 75.950 ;
        RECT 99.960 74.720 100.130 75.720 ;
        RECT 101.510 74.720 101.680 75.720 ;
        RECT 100.300 74.490 101.340 74.660 ;
        RECT 99.960 73.430 100.130 74.430 ;
        RECT 101.510 73.430 101.680 74.430 ;
        RECT 100.300 73.200 101.340 73.370 ;
        RECT 99.450 72.800 99.620 73.050 ;
        RECT 102.020 72.800 102.190 77.640 ;
        RECT 99.450 72.630 102.190 72.800 ;
        RECT 113.620 71.480 113.860 78.840 ;
        RECT 114.540 78.520 115.580 78.690 ;
        RECT 114.200 76.460 114.370 78.460 ;
        RECT 115.750 76.460 115.920 78.460 ;
        RECT 114.540 76.230 115.580 76.400 ;
        RECT 114.200 74.170 114.370 76.170 ;
        RECT 115.750 74.170 115.920 76.170 ;
        RECT 114.540 73.940 115.580 74.110 ;
        RECT 114.200 71.880 114.370 73.880 ;
        RECT 115.750 71.880 115.920 73.880 ;
        RECT 114.540 71.650 115.580 71.820 ;
        RECT 113.690 71.250 113.860 71.480 ;
        RECT 116.260 71.250 116.430 79.090 ;
        RECT 122.520 78.260 126.020 78.430 ;
        RECT 122.520 75.370 122.690 78.260 ;
        RECT 125.850 78.000 126.020 78.260 ;
        RECT 123.415 77.690 125.125 77.860 ;
        RECT 123.030 77.280 123.200 77.630 ;
        RECT 125.340 77.280 125.510 77.630 ;
        RECT 123.415 77.050 125.125 77.220 ;
        RECT 123.030 76.640 123.200 76.990 ;
        RECT 125.340 76.640 125.510 76.990 ;
        RECT 123.415 76.410 125.125 76.580 ;
        RECT 123.030 76.000 123.200 76.350 ;
        RECT 125.340 76.000 125.510 76.350 ;
        RECT 123.415 75.770 125.125 75.940 ;
        RECT 125.850 75.630 126.100 78.000 ;
        RECT 125.850 75.370 126.020 75.630 ;
        RECT 122.520 75.200 126.020 75.370 ;
        RECT 113.690 71.080 116.430 71.250 ;
        RECT 122.320 69.700 126.150 69.870 ;
        RECT 105.220 64.220 107.960 64.390 ;
        RECT 105.220 63.990 105.390 64.220 ;
        RECT 104.990 63.040 105.390 63.990 ;
        RECT 105.730 63.350 105.900 63.680 ;
        RECT 106.070 63.650 107.110 63.820 ;
        RECT 106.070 63.210 107.110 63.380 ;
        RECT 107.280 63.350 107.450 63.680 ;
        RECT 105.220 62.810 105.390 63.040 ;
        RECT 107.790 62.810 107.960 64.220 ;
        RECT 105.220 62.640 107.960 62.810 ;
        RECT 110.550 64.270 114.380 64.440 ;
        RECT 110.550 62.660 110.720 64.270 ;
        RECT 114.210 64.030 114.380 64.270 ;
        RECT 111.445 63.700 113.485 63.870 ;
        RECT 111.060 63.290 111.230 63.640 ;
        RECT 113.700 63.290 113.870 63.640 ;
        RECT 111.445 63.060 113.485 63.230 ;
        RECT 114.210 62.920 114.480 64.030 ;
        RECT 114.210 62.660 114.380 62.920 ;
        RECT 110.550 62.490 114.380 62.660 ;
        RECT 110.550 60.130 114.380 60.300 ;
        RECT 105.220 59.540 108.460 59.710 ;
        RECT 105.220 59.300 105.390 59.540 ;
        RECT 104.970 57.850 105.390 59.300 ;
        RECT 105.730 58.650 105.900 58.980 ;
        RECT 106.070 58.970 107.610 59.140 ;
        RECT 106.070 58.490 107.610 58.660 ;
        RECT 106.070 58.010 107.610 58.180 ;
        RECT 107.780 58.170 107.950 58.500 ;
        RECT 105.220 57.610 105.390 57.850 ;
        RECT 108.290 57.610 108.460 59.540 ;
        RECT 105.220 57.440 108.460 57.610 ;
        RECT 110.550 57.240 110.720 60.130 ;
        RECT 114.210 59.880 114.380 60.130 ;
        RECT 111.445 59.560 113.485 59.730 ;
        RECT 111.060 59.150 111.230 59.500 ;
        RECT 113.700 59.150 113.870 59.500 ;
        RECT 111.445 58.920 113.485 59.090 ;
        RECT 111.060 58.510 111.230 58.860 ;
        RECT 113.700 58.510 113.870 58.860 ;
        RECT 111.445 58.280 113.485 58.450 ;
        RECT 111.060 57.870 111.230 58.220 ;
        RECT 113.700 57.870 113.870 58.220 ;
        RECT 111.445 57.640 113.485 57.810 ;
        RECT 114.210 57.480 114.450 59.880 ;
        RECT 114.210 57.240 114.380 57.480 ;
        RECT 110.550 57.070 114.380 57.240 ;
        RECT 110.550 53.910 115.380 54.080 ;
        RECT 103.780 52.710 108.520 52.880 ;
        RECT 103.780 52.450 103.950 52.710 ;
        RECT 103.460 50.550 103.950 52.450 ;
        RECT 104.290 51.820 104.460 52.150 ;
        RECT 104.630 52.140 107.670 52.310 ;
        RECT 104.630 51.660 107.670 51.830 ;
        RECT 104.290 50.860 104.460 51.190 ;
        RECT 104.630 51.180 107.670 51.350 ;
        RECT 107.840 51.340 108.010 51.670 ;
        RECT 104.630 50.700 107.670 50.870 ;
        RECT 103.780 50.300 103.950 50.550 ;
        RECT 108.350 50.300 108.520 52.710 ;
        RECT 103.780 50.130 108.520 50.300 ;
        RECT 110.550 49.100 110.720 53.910 ;
        RECT 115.210 53.650 115.380 53.910 ;
        RECT 111.445 53.340 114.485 53.510 ;
        RECT 111.060 52.930 111.230 53.280 ;
        RECT 114.700 52.930 114.870 53.280 ;
        RECT 111.445 52.700 114.485 52.870 ;
        RECT 111.060 52.290 111.230 52.640 ;
        RECT 114.700 52.290 114.870 52.640 ;
        RECT 111.445 52.060 114.485 52.230 ;
        RECT 111.060 51.650 111.230 52.000 ;
        RECT 114.700 51.650 114.870 52.000 ;
        RECT 111.445 51.420 114.485 51.590 ;
        RECT 111.060 51.010 111.230 51.360 ;
        RECT 114.700 51.010 114.870 51.360 ;
        RECT 111.445 50.780 114.485 50.950 ;
        RECT 111.060 50.370 111.230 50.720 ;
        RECT 114.700 50.370 114.870 50.720 ;
        RECT 111.445 50.140 114.485 50.310 ;
        RECT 111.060 49.730 111.230 50.080 ;
        RECT 114.700 49.730 114.870 50.080 ;
        RECT 111.445 49.500 114.485 49.670 ;
        RECT 115.210 49.370 115.440 53.650 ;
        RECT 115.210 49.100 115.380 49.370 ;
        RECT 110.550 48.930 115.380 49.100 ;
        RECT 122.320 48.990 122.490 69.700 ;
        RECT 125.980 69.430 126.150 69.700 ;
        RECT 123.215 69.130 125.255 69.300 ;
        RECT 122.830 66.070 123.000 69.070 ;
        RECT 125.470 66.070 125.640 69.070 ;
        RECT 123.215 65.840 125.255 66.010 ;
        RECT 122.830 62.780 123.000 65.780 ;
        RECT 125.470 62.780 125.640 65.780 ;
        RECT 123.215 62.550 125.255 62.720 ;
        RECT 122.830 59.490 123.000 62.490 ;
        RECT 125.470 59.490 125.640 62.490 ;
        RECT 123.215 59.260 125.255 59.430 ;
        RECT 122.830 56.200 123.000 59.200 ;
        RECT 125.470 56.200 125.640 59.200 ;
        RECT 123.215 55.970 125.255 56.140 ;
        RECT 122.830 52.910 123.000 55.910 ;
        RECT 125.470 52.910 125.640 55.910 ;
        RECT 123.215 52.680 125.255 52.850 ;
        RECT 122.830 49.620 123.000 52.620 ;
        RECT 125.470 49.620 125.640 52.620 ;
        RECT 123.215 49.390 125.255 49.560 ;
        RECT 125.980 49.250 126.230 69.430 ;
        RECT 125.980 48.990 126.150 49.250 ;
        RECT 122.320 48.820 126.150 48.990 ;
      LAYER mcon ;
        RECT 96.720 136.960 99.600 137.130 ;
        RECT 96.300 133.980 96.470 136.820 ;
        RECT 99.850 133.980 100.020 136.820 ;
        RECT 96.720 133.670 99.600 133.840 ;
        RECT 105.900 137.530 109.750 137.750 ;
        RECT 106.380 136.960 109.260 137.130 ;
        RECT 105.960 136.720 106.130 136.890 ;
        RECT 106.380 136.480 109.260 136.650 ;
        RECT 109.510 136.240 109.680 136.410 ;
        RECT 106.380 136.000 109.260 136.170 ;
        RECT 105.960 135.760 106.130 135.930 ;
        RECT 106.380 135.520 109.260 135.690 ;
        RECT 109.510 135.280 109.680 135.450 ;
        RECT 106.380 135.040 109.260 135.210 ;
        RECT 105.960 134.800 106.130 134.970 ;
        RECT 106.380 134.560 109.260 134.730 ;
        RECT 109.510 134.320 109.680 134.490 ;
        RECT 106.380 134.080 109.260 134.250 ;
        RECT 105.960 133.840 106.130 134.010 ;
        RECT 106.380 133.600 109.260 133.770 ;
        RECT 115.040 137.530 118.940 137.730 ;
        RECT 115.555 136.960 118.435 137.130 ;
        RECT 115.090 136.630 115.260 136.820 ;
        RECT 118.730 136.630 118.900 136.820 ;
        RECT 115.555 136.320 118.435 136.490 ;
        RECT 115.090 135.990 115.260 136.180 ;
        RECT 118.730 135.990 118.900 136.180 ;
        RECT 115.555 135.680 118.435 135.850 ;
        RECT 115.090 135.350 115.260 135.540 ;
        RECT 118.730 135.350 118.900 135.540 ;
        RECT 115.555 135.040 118.435 135.210 ;
        RECT 115.090 134.710 115.260 134.900 ;
        RECT 118.730 134.710 118.900 134.900 ;
        RECT 115.555 134.400 118.435 134.570 ;
        RECT 115.090 134.070 115.260 134.260 ;
        RECT 118.730 134.070 118.900 134.260 ;
        RECT 115.555 133.760 118.435 133.930 ;
        RECT 115.090 133.430 115.260 133.620 ;
        RECT 118.730 133.430 118.900 133.620 ;
        RECT 115.555 133.120 118.435 133.290 ;
        RECT 115.090 132.790 115.260 132.980 ;
        RECT 118.730 132.790 118.900 132.980 ;
        RECT 115.555 132.480 118.435 132.650 ;
        RECT 123.945 136.850 126.825 137.020 ;
        RECT 123.480 133.870 123.650 136.710 ;
        RECT 127.120 133.870 127.290 136.710 ;
        RECT 123.945 133.560 126.825 133.730 ;
        RECT 97.300 121.790 101.180 121.960 ;
        RECT 96.880 118.810 97.050 121.650 ;
        RECT 101.430 118.810 101.600 121.650 ;
        RECT 97.300 118.500 101.180 118.670 ;
        RECT 96.880 115.520 97.050 118.360 ;
        RECT 101.430 115.520 101.600 118.360 ;
        RECT 97.300 115.210 101.180 115.380 ;
        RECT 96.880 112.230 97.050 115.070 ;
        RECT 101.430 112.230 101.600 115.070 ;
        RECT 97.300 111.920 101.180 112.090 ;
        RECT 97.360 106.190 101.240 106.360 ;
        RECT 96.940 103.210 97.110 106.050 ;
        RECT 101.490 103.210 101.660 106.050 ;
        RECT 97.360 102.900 101.240 103.070 ;
        RECT 96.940 99.920 97.110 102.760 ;
        RECT 101.490 99.920 101.660 102.760 ;
        RECT 97.360 99.610 101.240 99.780 ;
        RECT 96.940 96.630 97.110 99.470 ;
        RECT 101.490 96.630 101.660 99.470 ;
        RECT 97.360 96.320 101.240 96.490 ;
        RECT 108.175 118.140 109.555 118.310 ;
        RECT 107.710 117.460 107.880 118.000 ;
        RECT 109.850 117.460 110.020 118.000 ;
        RECT 108.175 117.150 109.555 117.320 ;
        RECT 107.710 116.470 107.880 117.010 ;
        RECT 109.850 116.470 110.020 117.010 ;
        RECT 108.175 116.160 109.555 116.330 ;
        RECT 107.710 115.480 107.880 116.020 ;
        RECT 109.850 115.480 110.020 116.020 ;
        RECT 108.175 115.170 109.555 115.340 ;
        RECT 107.710 114.490 107.880 115.030 ;
        RECT 109.850 114.490 110.020 115.030 ;
        RECT 108.175 114.180 109.555 114.350 ;
        RECT 107.710 113.500 107.880 114.040 ;
        RECT 109.850 113.500 110.020 114.040 ;
        RECT 108.175 113.190 109.555 113.360 ;
        RECT 107.710 112.510 107.880 113.050 ;
        RECT 109.850 112.510 110.020 113.050 ;
        RECT 108.175 112.200 109.555 112.370 ;
        RECT 107.710 111.520 107.880 112.060 ;
        RECT 109.850 111.520 110.020 112.060 ;
        RECT 108.175 111.210 109.555 111.380 ;
        RECT 107.710 110.530 107.880 111.070 ;
        RECT 109.850 110.530 110.020 111.070 ;
        RECT 108.175 110.220 109.555 110.390 ;
        RECT 107.710 109.540 107.880 110.080 ;
        RECT 109.850 109.540 110.020 110.080 ;
        RECT 108.175 109.230 109.555 109.400 ;
        RECT 107.710 108.550 107.880 109.090 ;
        RECT 109.850 108.550 110.020 109.090 ;
        RECT 108.175 108.240 109.555 108.410 ;
        RECT 107.710 107.560 107.880 108.100 ;
        RECT 109.850 107.560 110.020 108.100 ;
        RECT 108.175 107.250 109.555 107.420 ;
        RECT 107.710 106.570 107.880 107.110 ;
        RECT 109.850 106.570 110.020 107.110 ;
        RECT 108.175 106.260 109.555 106.430 ;
        RECT 107.710 105.580 107.880 106.120 ;
        RECT 109.850 105.580 110.020 106.120 ;
        RECT 108.175 105.270 109.555 105.440 ;
        RECT 107.710 104.590 107.880 105.130 ;
        RECT 109.850 104.590 110.020 105.130 ;
        RECT 108.175 104.280 109.555 104.450 ;
        RECT 107.710 103.600 107.880 104.140 ;
        RECT 109.850 103.600 110.020 104.140 ;
        RECT 108.175 103.290 109.555 103.460 ;
        RECT 107.710 102.610 107.880 103.150 ;
        RECT 109.850 102.610 110.020 103.150 ;
        RECT 108.175 102.300 109.555 102.470 ;
        RECT 107.710 101.620 107.880 102.160 ;
        RECT 109.850 101.620 110.020 102.160 ;
        RECT 108.175 101.310 109.555 101.480 ;
        RECT 107.710 100.630 107.880 101.170 ;
        RECT 109.850 100.630 110.020 101.170 ;
        RECT 108.175 100.320 109.555 100.490 ;
        RECT 116.005 118.140 117.385 118.310 ;
        RECT 115.540 117.460 115.710 118.000 ;
        RECT 117.680 117.460 117.850 118.000 ;
        RECT 116.005 117.150 117.385 117.320 ;
        RECT 115.540 116.470 115.710 117.010 ;
        RECT 117.680 116.470 117.850 117.010 ;
        RECT 116.005 116.160 117.385 116.330 ;
        RECT 115.540 115.480 115.710 116.020 ;
        RECT 117.680 115.480 117.850 116.020 ;
        RECT 116.005 115.170 117.385 115.340 ;
        RECT 115.540 114.490 115.710 115.030 ;
        RECT 117.680 114.490 117.850 115.030 ;
        RECT 116.005 114.180 117.385 114.350 ;
        RECT 115.540 113.500 115.710 114.040 ;
        RECT 117.680 113.500 117.850 114.040 ;
        RECT 116.005 113.190 117.385 113.360 ;
        RECT 115.540 112.510 115.710 113.050 ;
        RECT 117.680 112.510 117.850 113.050 ;
        RECT 116.005 112.200 117.385 112.370 ;
        RECT 115.540 111.520 115.710 112.060 ;
        RECT 117.680 111.520 117.850 112.060 ;
        RECT 116.005 111.210 117.385 111.380 ;
        RECT 115.540 110.530 115.710 111.070 ;
        RECT 117.680 110.530 117.850 111.070 ;
        RECT 116.005 110.220 117.385 110.390 ;
        RECT 115.540 109.540 115.710 110.080 ;
        RECT 117.680 109.540 117.850 110.080 ;
        RECT 116.005 109.230 117.385 109.400 ;
        RECT 115.540 108.550 115.710 109.090 ;
        RECT 117.680 108.550 117.850 109.090 ;
        RECT 116.005 108.240 117.385 108.410 ;
        RECT 115.540 107.560 115.710 108.100 ;
        RECT 117.680 107.560 117.850 108.100 ;
        RECT 116.005 107.250 117.385 107.420 ;
        RECT 115.540 106.570 115.710 107.110 ;
        RECT 117.680 106.570 117.850 107.110 ;
        RECT 116.005 106.260 117.385 106.430 ;
        RECT 115.540 105.580 115.710 106.120 ;
        RECT 117.680 105.580 117.850 106.120 ;
        RECT 116.005 105.270 117.385 105.440 ;
        RECT 115.540 104.590 115.710 105.130 ;
        RECT 117.680 104.590 117.850 105.130 ;
        RECT 116.005 104.280 117.385 104.450 ;
        RECT 115.540 103.600 115.710 104.140 ;
        RECT 117.680 103.600 117.850 104.140 ;
        RECT 116.005 103.290 117.385 103.460 ;
        RECT 115.540 102.610 115.710 103.150 ;
        RECT 117.680 102.610 117.850 103.150 ;
        RECT 116.005 102.300 117.385 102.470 ;
        RECT 115.540 101.620 115.710 102.160 ;
        RECT 117.680 101.620 117.850 102.160 ;
        RECT 116.005 101.310 117.385 101.480 ;
        RECT 115.540 100.630 115.710 101.170 ;
        RECT 117.680 100.630 117.850 101.170 ;
        RECT 116.005 100.320 117.385 100.490 ;
        RECT 100.350 91.040 101.230 91.210 ;
        RECT 99.930 90.060 100.100 90.900 ;
        RECT 101.480 90.060 101.650 90.900 ;
        RECT 100.350 89.750 101.230 89.920 ;
        RECT 99.930 88.770 100.100 89.610 ;
        RECT 101.480 88.770 101.650 89.610 ;
        RECT 100.350 88.460 101.230 88.630 ;
        RECT 99.930 87.480 100.100 88.320 ;
        RECT 101.480 87.480 101.650 88.320 ;
        RECT 100.350 87.170 101.230 87.340 ;
        RECT 113.535 91.550 115.555 91.720 ;
        RECT 113.070 91.220 113.240 91.410 ;
        RECT 115.850 91.220 116.020 91.410 ;
        RECT 113.535 90.910 115.555 91.080 ;
        RECT 113.070 90.580 113.240 90.770 ;
        RECT 115.850 90.580 116.020 90.770 ;
        RECT 113.535 90.270 115.555 90.440 ;
        RECT 113.070 89.940 113.240 90.130 ;
        RECT 115.850 89.940 116.020 90.130 ;
        RECT 113.535 89.630 115.555 89.800 ;
        RECT 113.070 89.300 113.240 89.490 ;
        RECT 115.850 89.300 116.020 89.490 ;
        RECT 113.535 88.990 115.555 89.160 ;
        RECT 113.070 88.660 113.240 88.850 ;
        RECT 115.850 88.660 116.020 88.850 ;
        RECT 113.535 88.350 115.555 88.520 ;
        RECT 113.070 88.020 113.240 88.210 ;
        RECT 115.850 88.020 116.020 88.210 ;
        RECT 113.535 87.710 115.555 87.880 ;
        RECT 113.070 87.380 113.240 87.570 ;
        RECT 115.850 87.380 116.020 87.570 ;
        RECT 113.535 87.070 115.555 87.240 ;
        RECT 123.845 114.770 125.725 114.940 ;
        RECT 123.380 111.790 123.550 114.630 ;
        RECT 126.020 111.790 126.190 114.630 ;
        RECT 123.845 111.480 125.725 111.650 ;
        RECT 123.380 108.500 123.550 111.340 ;
        RECT 126.020 108.500 126.190 111.340 ;
        RECT 123.845 108.190 125.725 108.360 ;
        RECT 123.380 105.210 123.550 108.050 ;
        RECT 126.020 105.210 126.190 108.050 ;
        RECT 123.845 104.900 125.725 105.070 ;
        RECT 123.380 101.920 123.550 104.760 ;
        RECT 126.020 101.920 126.190 104.760 ;
        RECT 123.845 101.610 125.725 101.780 ;
        RECT 123.380 98.630 123.550 101.470 ;
        RECT 126.020 98.630 126.190 101.470 ;
        RECT 123.845 98.320 125.725 98.490 ;
        RECT 123.380 95.340 123.550 98.180 ;
        RECT 126.020 95.340 126.190 98.180 ;
        RECT 123.845 95.030 125.725 95.200 ;
        RECT 123.380 92.050 123.550 94.890 ;
        RECT 126.020 92.050 126.190 94.890 ;
        RECT 123.845 91.740 125.725 91.910 ;
        RECT 123.380 88.760 123.550 91.600 ;
        RECT 126.020 88.760 126.190 91.600 ;
        RECT 123.845 88.450 125.725 88.620 ;
        RECT 123.380 85.470 123.550 88.310 ;
        RECT 126.020 85.470 126.190 88.310 ;
        RECT 123.845 85.160 125.725 85.330 ;
        RECT 100.380 77.070 101.260 77.240 ;
        RECT 99.960 76.090 100.130 76.930 ;
        RECT 101.510 76.090 101.680 76.930 ;
        RECT 100.380 75.780 101.260 75.950 ;
        RECT 99.960 74.800 100.130 75.640 ;
        RECT 101.510 74.800 101.680 75.640 ;
        RECT 100.380 74.490 101.260 74.660 ;
        RECT 99.960 73.510 100.130 74.350 ;
        RECT 101.510 73.510 101.680 74.350 ;
        RECT 100.380 73.200 101.260 73.370 ;
        RECT 114.620 78.520 115.500 78.690 ;
        RECT 114.200 76.540 114.370 78.380 ;
        RECT 115.750 76.540 115.920 78.380 ;
        RECT 114.620 76.230 115.500 76.400 ;
        RECT 114.200 74.250 114.370 76.090 ;
        RECT 115.750 74.250 115.920 76.090 ;
        RECT 114.620 73.940 115.500 74.110 ;
        RECT 114.200 71.960 114.370 73.800 ;
        RECT 115.750 71.960 115.920 73.800 ;
        RECT 114.620 71.650 115.500 71.820 ;
        RECT 123.495 77.690 125.045 77.860 ;
        RECT 123.030 77.360 123.200 77.550 ;
        RECT 125.340 77.360 125.510 77.550 ;
        RECT 123.495 77.050 125.045 77.220 ;
        RECT 123.030 76.720 123.200 76.910 ;
        RECT 125.340 76.720 125.510 76.910 ;
        RECT 123.495 76.410 125.045 76.580 ;
        RECT 123.030 76.080 123.200 76.270 ;
        RECT 125.340 76.080 125.510 76.270 ;
        RECT 123.495 75.770 125.045 75.940 ;
        RECT 106.150 63.650 107.030 63.820 ;
        RECT 105.730 63.430 105.900 63.600 ;
        RECT 107.280 63.430 107.450 63.600 ;
        RECT 106.150 63.210 107.030 63.380 ;
        RECT 111.525 63.700 113.405 63.870 ;
        RECT 111.060 63.370 111.230 63.560 ;
        RECT 113.700 63.370 113.870 63.560 ;
        RECT 111.525 63.060 113.405 63.230 ;
        RECT 106.150 58.970 107.530 59.140 ;
        RECT 105.730 58.730 105.900 58.900 ;
        RECT 106.150 58.490 107.530 58.660 ;
        RECT 107.780 58.250 107.950 58.420 ;
        RECT 106.150 58.010 107.530 58.180 ;
        RECT 111.525 59.560 113.405 59.730 ;
        RECT 111.060 59.230 111.230 59.420 ;
        RECT 113.700 59.230 113.870 59.420 ;
        RECT 111.525 58.920 113.405 59.090 ;
        RECT 111.060 58.590 111.230 58.780 ;
        RECT 113.700 58.590 113.870 58.780 ;
        RECT 111.525 58.280 113.405 58.450 ;
        RECT 111.060 57.950 111.230 58.140 ;
        RECT 113.700 57.950 113.870 58.140 ;
        RECT 111.525 57.640 113.405 57.810 ;
        RECT 104.710 52.140 107.590 52.310 ;
        RECT 104.290 51.900 104.460 52.070 ;
        RECT 104.710 51.660 107.590 51.830 ;
        RECT 107.840 51.420 108.010 51.590 ;
        RECT 104.710 51.180 107.590 51.350 ;
        RECT 104.290 50.940 104.460 51.110 ;
        RECT 104.710 50.700 107.590 50.870 ;
        RECT 111.525 53.340 114.405 53.510 ;
        RECT 111.060 53.010 111.230 53.200 ;
        RECT 114.700 53.010 114.870 53.200 ;
        RECT 111.525 52.700 114.405 52.870 ;
        RECT 111.060 52.370 111.230 52.560 ;
        RECT 114.700 52.370 114.870 52.560 ;
        RECT 111.525 52.060 114.405 52.230 ;
        RECT 111.060 51.730 111.230 51.920 ;
        RECT 114.700 51.730 114.870 51.920 ;
        RECT 111.525 51.420 114.405 51.590 ;
        RECT 111.060 51.090 111.230 51.280 ;
        RECT 114.700 51.090 114.870 51.280 ;
        RECT 111.525 50.780 114.405 50.950 ;
        RECT 111.060 50.450 111.230 50.640 ;
        RECT 114.700 50.450 114.870 50.640 ;
        RECT 111.525 50.140 114.405 50.310 ;
        RECT 111.060 49.810 111.230 50.000 ;
        RECT 114.700 49.810 114.870 50.000 ;
        RECT 111.525 49.500 114.405 49.670 ;
        RECT 123.295 69.130 125.175 69.300 ;
        RECT 122.830 66.150 123.000 68.990 ;
        RECT 125.470 66.150 125.640 68.990 ;
        RECT 123.295 65.840 125.175 66.010 ;
        RECT 122.830 62.860 123.000 65.700 ;
        RECT 125.470 62.860 125.640 65.700 ;
        RECT 123.295 62.550 125.175 62.720 ;
        RECT 122.830 59.570 123.000 62.410 ;
        RECT 125.470 59.570 125.640 62.410 ;
        RECT 123.295 59.260 125.175 59.430 ;
        RECT 122.830 56.280 123.000 59.120 ;
        RECT 125.470 56.280 125.640 59.120 ;
        RECT 123.295 55.970 125.175 56.140 ;
        RECT 122.830 52.990 123.000 55.830 ;
        RECT 125.470 52.990 125.640 55.830 ;
        RECT 123.295 52.680 125.175 52.850 ;
        RECT 122.830 49.700 123.000 52.540 ;
        RECT 125.470 49.700 125.640 52.540 ;
        RECT 123.295 49.390 125.175 49.560 ;
        RECT 125.990 49.250 126.230 69.430 ;
      LAYER met1 ;
        RECT 90.710 153.455 93.855 153.675 ;
        RECT 87.485 150.745 93.855 153.455 ;
        RECT 90.710 142.280 93.855 150.745 ;
        RECT 118.920 147.490 120.300 147.520 ;
        RECT 111.930 146.110 120.300 147.490 ;
        RECT 111.930 142.630 113.310 146.110 ;
        RECT 118.920 146.080 120.300 146.110 ;
        RECT 90.530 142.270 94.550 142.280 ;
        RECT 90.530 139.990 110.030 142.270 ;
        RECT 90.530 139.910 110.040 139.990 ;
        RECT 90.530 137.510 94.550 139.910 ;
        RECT 90.530 133.270 95.990 137.510 ;
        RECT 96.700 137.160 99.630 139.910 ;
        RECT 105.710 137.500 110.040 139.910 ;
        RECT 108.830 137.160 109.320 137.220 ;
        RECT 96.660 136.930 99.660 137.160 ;
        RECT 90.530 122.140 94.550 133.270 ;
        RECT 96.270 130.710 96.510 136.900 ;
        RECT 96.730 133.870 99.630 133.890 ;
        RECT 96.660 133.640 99.660 133.870 ;
        RECT 96.730 133.470 99.630 133.640 ;
        RECT 97.380 132.640 98.220 133.470 ;
        RECT 97.385 130.710 98.215 132.640 ;
        RECT 99.810 130.710 100.110 136.910 ;
        RECT 103.460 131.920 104.080 132.480 ;
        RECT 103.490 130.710 104.050 131.920 ;
        RECT 96.270 130.110 104.050 130.710 ;
        RECT 105.810 130.670 106.160 136.980 ;
        RECT 106.320 136.930 109.320 137.160 ;
        RECT 108.830 136.830 109.320 136.930 ;
        RECT 106.390 136.680 106.880 136.760 ;
        RECT 106.320 136.450 109.320 136.680 ;
        RECT 106.390 136.370 106.880 136.450 ;
        RECT 108.830 136.200 109.320 136.280 ;
        RECT 106.320 135.970 109.320 136.200 ;
        RECT 108.830 135.890 109.320 135.970 ;
        RECT 106.390 135.720 106.880 135.800 ;
        RECT 106.320 135.490 109.320 135.720 ;
        RECT 106.390 135.410 106.880 135.490 ;
        RECT 108.830 135.240 109.320 135.320 ;
        RECT 106.320 135.010 109.320 135.240 ;
        RECT 108.830 134.930 109.320 135.010 ;
        RECT 106.390 134.760 106.880 134.840 ;
        RECT 106.320 134.530 109.320 134.760 ;
        RECT 106.390 134.450 106.880 134.530 ;
        RECT 108.830 134.280 109.320 134.360 ;
        RECT 106.320 134.050 109.320 134.280 ;
        RECT 108.830 133.970 109.320 134.050 ;
        RECT 106.390 133.800 106.880 133.880 ;
        RECT 106.320 133.570 109.320 133.800 ;
        RECT 106.390 133.490 106.880 133.570 ;
        RECT 108.015 130.670 108.585 132.570 ;
        RECT 109.460 130.670 109.810 136.530 ;
        RECT 111.750 133.380 113.315 142.630 ;
        RECT 129.020 142.420 131.975 162.360 ;
        RECT 114.970 140.130 132.620 142.420 ;
        RECT 114.960 140.060 132.620 140.130 ;
        RECT 114.960 137.460 118.980 140.060 ;
        RECT 115.570 137.160 116.050 137.170 ;
        RECT 114.990 131.290 115.300 136.960 ;
        RECT 115.495 136.930 118.495 137.160 ;
        RECT 124.080 137.050 126.610 140.060 ;
        RECT 128.600 137.590 132.620 140.060 ;
        RECT 115.570 136.790 116.050 136.930 ;
        RECT 117.970 136.520 118.450 136.600 ;
        RECT 115.495 136.290 118.495 136.520 ;
        RECT 117.970 136.220 118.450 136.290 ;
        RECT 115.550 135.880 116.030 135.950 ;
        RECT 115.495 135.650 118.495 135.880 ;
        RECT 115.550 135.570 116.030 135.650 ;
        RECT 117.970 135.240 118.450 135.310 ;
        RECT 115.495 135.010 118.495 135.240 ;
        RECT 117.970 134.930 118.450 135.010 ;
        RECT 115.550 134.600 116.030 134.680 ;
        RECT 115.495 134.370 118.495 134.600 ;
        RECT 115.550 134.300 116.030 134.370 ;
        RECT 117.970 133.960 118.450 134.040 ;
        RECT 115.495 133.730 118.495 133.960 ;
        RECT 117.970 133.660 118.450 133.730 ;
        RECT 115.550 133.320 116.030 133.390 ;
        RECT 115.495 133.090 118.495 133.320 ;
        RECT 115.550 133.010 116.030 133.090 ;
        RECT 117.970 132.680 118.450 132.760 ;
        RECT 115.495 132.450 118.495 132.680 ;
        RECT 117.970 132.380 118.450 132.450 ;
        RECT 114.990 130.710 116.130 131.290 ;
        RECT 114.990 130.670 116.100 130.710 ;
        RECT 105.800 130.400 116.100 130.670 ;
        RECT 118.650 130.400 118.960 136.960 ;
        RECT 123.410 136.770 123.660 136.850 ;
        RECT 123.885 136.820 126.885 137.050 ;
        RECT 127.060 136.770 127.310 136.850 ;
        RECT 123.410 133.810 123.680 136.770 ;
        RECT 127.060 133.810 127.320 136.770 ;
        RECT 123.410 132.160 123.660 133.810 ;
        RECT 123.885 133.530 126.885 133.760 ;
        RECT 125.030 132.160 126.180 133.530 ;
        RECT 127.060 132.160 127.310 133.810 ;
        RECT 127.600 132.970 132.620 137.590 ;
        RECT 123.410 131.985 127.310 132.160 ;
        RECT 121.315 131.435 127.315 131.985 ;
        RECT 120.440 131.250 120.980 131.280 ;
        RECT 121.315 131.250 121.865 131.435 ;
        RECT 120.440 130.710 121.865 131.250 ;
        RECT 120.440 130.680 120.980 130.710 ;
        RECT 121.315 130.705 121.865 130.710 ;
        RECT 96.270 130.030 104.030 130.110 ;
        RECT 105.800 130.090 118.965 130.400 ;
        RECT 105.800 130.070 115.440 130.090 ;
        RECT 100.800 127.520 101.730 130.030 ;
        RECT 125.630 128.345 126.220 131.435 ;
        RECT 125.600 127.755 126.250 128.345 ;
        RECT 100.800 126.580 104.730 127.520 ;
        RECT 100.800 125.510 101.730 126.580 ;
        RECT 96.850 124.070 101.740 125.510 ;
        RECT 90.530 111.700 96.570 122.140 ;
        RECT 96.850 112.140 97.100 124.070 ;
        RECT 100.540 121.990 101.170 122.080 ;
        RECT 97.240 121.760 101.240 121.990 ;
        RECT 100.540 121.660 101.170 121.760 ;
        RECT 97.310 118.700 97.940 118.810 ;
        RECT 97.240 118.470 101.240 118.700 ;
        RECT 97.310 118.390 97.940 118.470 ;
        RECT 100.540 115.410 101.170 115.500 ;
        RECT 97.240 115.180 101.240 115.410 ;
        RECT 100.540 115.080 101.170 115.180 ;
        RECT 97.310 112.120 97.940 112.200 ;
        RECT 97.240 111.890 101.240 112.120 ;
        RECT 101.400 111.940 101.740 124.070 ;
        RECT 97.310 111.780 97.940 111.890 ;
        RECT 90.530 110.520 94.550 111.700 ;
        RECT 90.530 109.770 98.040 110.520 ;
        RECT 90.530 106.690 94.550 109.770 ;
        RECT 101.450 108.410 101.830 108.420 ;
        RECT 103.790 108.410 104.730 126.580 ;
        RECT 110.770 123.460 112.160 123.465 ;
        RECT 118.480 123.460 120.070 123.465 ;
        RECT 128.600 123.460 132.620 132.970 ;
        RECT 110.770 120.240 132.620 123.460 ;
        RECT 110.770 118.560 112.160 120.240 ;
        RECT 109.150 118.340 109.560 118.420 ;
        RECT 96.910 107.470 104.730 108.410 ;
        RECT 90.530 96.090 96.630 106.690 ;
        RECT 96.910 96.570 97.160 107.470 ;
        RECT 100.540 106.390 101.250 106.500 ;
        RECT 97.300 106.160 101.300 106.390 ;
        RECT 100.540 106.030 101.250 106.160 ;
        RECT 97.360 103.100 98.070 103.210 ;
        RECT 97.300 102.870 101.300 103.100 ;
        RECT 97.360 102.740 98.070 102.870 ;
        RECT 100.540 99.810 101.250 99.930 ;
        RECT 97.300 99.580 101.300 99.810 ;
        RECT 100.540 99.460 101.250 99.580 ;
        RECT 97.360 96.520 98.070 96.640 ;
        RECT 97.300 96.290 101.300 96.520 ;
        RECT 101.450 96.450 101.830 107.470 ;
        RECT 107.610 98.650 107.930 118.140 ;
        RECT 108.115 118.110 109.615 118.340 ;
        RECT 109.150 118.030 109.560 118.110 ;
        RECT 108.170 117.350 108.580 117.430 ;
        RECT 108.115 117.120 109.615 117.350 ;
        RECT 108.170 117.040 108.580 117.120 ;
        RECT 109.150 116.360 109.560 116.440 ;
        RECT 108.115 116.130 109.615 116.360 ;
        RECT 109.150 116.050 109.560 116.130 ;
        RECT 108.170 115.370 108.580 115.450 ;
        RECT 108.115 115.140 109.615 115.370 ;
        RECT 108.170 115.060 108.580 115.140 ;
        RECT 109.150 114.380 109.560 114.460 ;
        RECT 108.115 114.150 109.615 114.380 ;
        RECT 109.150 114.070 109.560 114.150 ;
        RECT 108.170 113.390 108.580 113.470 ;
        RECT 108.115 113.160 109.615 113.390 ;
        RECT 108.170 113.080 108.580 113.160 ;
        RECT 109.150 112.400 109.560 112.480 ;
        RECT 108.115 112.170 109.615 112.400 ;
        RECT 109.150 112.090 109.560 112.170 ;
        RECT 108.170 111.410 108.580 111.500 ;
        RECT 108.115 111.180 109.615 111.410 ;
        RECT 108.170 111.110 108.580 111.180 ;
        RECT 109.150 110.420 109.560 110.500 ;
        RECT 108.115 110.190 109.615 110.420 ;
        RECT 109.150 110.110 109.560 110.190 ;
        RECT 108.170 109.430 108.580 109.520 ;
        RECT 108.115 109.200 109.615 109.430 ;
        RECT 108.170 109.130 108.580 109.200 ;
        RECT 109.150 108.440 109.560 108.520 ;
        RECT 108.115 108.210 109.615 108.440 ;
        RECT 109.150 108.130 109.560 108.210 ;
        RECT 108.170 107.450 108.580 107.530 ;
        RECT 108.115 107.220 109.615 107.450 ;
        RECT 108.170 107.140 108.580 107.220 ;
        RECT 109.150 106.460 109.560 106.540 ;
        RECT 108.115 106.230 109.615 106.460 ;
        RECT 109.150 106.150 109.560 106.230 ;
        RECT 108.170 105.470 108.580 105.560 ;
        RECT 108.115 105.240 109.615 105.470 ;
        RECT 108.170 105.170 108.580 105.240 ;
        RECT 109.150 104.480 109.560 104.560 ;
        RECT 108.115 104.250 109.615 104.480 ;
        RECT 109.150 104.170 109.560 104.250 ;
        RECT 108.170 103.490 108.580 103.570 ;
        RECT 108.115 103.260 109.615 103.490 ;
        RECT 108.170 103.180 108.580 103.260 ;
        RECT 109.150 102.500 109.560 102.580 ;
        RECT 108.115 102.270 109.615 102.500 ;
        RECT 109.150 102.190 109.560 102.270 ;
        RECT 108.170 101.510 108.580 101.590 ;
        RECT 108.115 101.280 109.615 101.510 ;
        RECT 108.170 101.200 108.580 101.280 ;
        RECT 109.150 100.520 109.560 100.600 ;
        RECT 108.115 100.290 109.615 100.520 ;
        RECT 109.150 100.210 109.560 100.290 ;
        RECT 109.770 98.650 110.090 118.140 ;
        RECT 110.300 100.010 112.160 118.560 ;
        RECT 118.480 118.440 120.070 120.240 ;
        RECT 116.940 118.340 117.470 118.420 ;
        RECT 115.945 118.110 117.470 118.340 ;
        RECT 115.430 98.650 115.750 118.080 ;
        RECT 116.940 118.030 117.470 118.110 ;
        RECT 115.980 117.350 116.510 117.430 ;
        RECT 115.945 117.120 117.445 117.350 ;
        RECT 115.980 117.040 116.510 117.120 ;
        RECT 116.940 116.360 117.470 116.440 ;
        RECT 115.945 116.130 117.470 116.360 ;
        RECT 116.940 116.050 117.470 116.130 ;
        RECT 115.980 115.370 116.510 115.460 ;
        RECT 115.945 115.140 117.445 115.370 ;
        RECT 115.980 115.070 116.510 115.140 ;
        RECT 116.940 114.380 117.470 114.460 ;
        RECT 115.945 114.150 117.470 114.380 ;
        RECT 116.940 114.070 117.470 114.150 ;
        RECT 115.980 113.390 116.510 113.480 ;
        RECT 115.945 113.160 117.445 113.390 ;
        RECT 115.980 113.090 116.510 113.160 ;
        RECT 116.940 112.400 117.470 112.490 ;
        RECT 115.945 112.170 117.470 112.400 ;
        RECT 116.940 112.100 117.470 112.170 ;
        RECT 115.980 111.410 116.510 111.490 ;
        RECT 115.945 111.180 117.445 111.410 ;
        RECT 115.980 111.100 116.510 111.180 ;
        RECT 116.940 110.420 117.470 110.510 ;
        RECT 115.945 110.190 117.470 110.420 ;
        RECT 116.940 110.120 117.470 110.190 ;
        RECT 115.980 109.430 116.510 109.510 ;
        RECT 115.945 109.200 117.445 109.430 ;
        RECT 115.980 109.120 116.510 109.200 ;
        RECT 116.940 108.440 117.470 108.520 ;
        RECT 115.945 108.210 117.470 108.440 ;
        RECT 116.940 108.130 117.470 108.210 ;
        RECT 115.980 107.450 116.510 107.540 ;
        RECT 115.945 107.220 117.445 107.450 ;
        RECT 115.980 107.150 116.510 107.220 ;
        RECT 116.940 106.460 117.470 106.540 ;
        RECT 115.945 106.230 117.470 106.460 ;
        RECT 116.940 106.150 117.470 106.230 ;
        RECT 115.980 105.470 116.510 105.560 ;
        RECT 115.945 105.240 117.445 105.470 ;
        RECT 115.980 105.170 116.510 105.240 ;
        RECT 116.940 104.480 117.470 104.570 ;
        RECT 115.945 104.250 117.470 104.480 ;
        RECT 116.940 104.180 117.470 104.250 ;
        RECT 115.980 103.490 116.510 103.580 ;
        RECT 115.945 103.260 117.445 103.490 ;
        RECT 115.980 103.190 116.510 103.260 ;
        RECT 116.940 102.500 117.470 102.580 ;
        RECT 115.945 102.270 117.470 102.500 ;
        RECT 116.940 102.190 117.470 102.270 ;
        RECT 115.980 101.510 116.510 101.600 ;
        RECT 115.945 101.280 117.445 101.510 ;
        RECT 115.980 101.210 116.510 101.280 ;
        RECT 116.940 100.520 117.470 100.600 ;
        RECT 115.945 100.290 117.470 100.520 ;
        RECT 116.940 100.210 117.470 100.290 ;
        RECT 117.640 98.650 117.960 118.100 ;
        RECT 118.110 100.910 120.070 118.440 ;
        RECT 125.630 116.930 126.220 117.985 ;
        RECT 123.350 116.340 126.220 116.930 ;
        RECT 118.110 100.150 120.090 100.910 ;
        RECT 107.590 98.185 117.970 98.650 ;
        RECT 106.435 97.590 117.970 98.185 ;
        RECT 106.435 97.560 111.070 97.590 ;
        RECT 106.435 97.495 111.065 97.560 ;
        RECT 97.360 96.170 98.070 96.290 ;
        RECT 90.530 94.590 94.550 96.090 ;
        RECT 106.435 95.755 107.125 97.495 ;
        RECT 90.530 93.790 98.150 94.590 ;
        RECT 90.530 91.430 94.550 93.790 ;
        RECT 113.010 93.710 113.680 95.135 ;
        RECT 113.010 93.040 116.070 93.710 ;
        RECT 100.340 92.680 100.700 92.710 ;
        RECT 98.700 92.320 100.700 92.680 ;
        RECT 98.700 91.430 99.060 92.320 ;
        RECT 100.340 92.290 100.700 92.320 ;
        RECT 90.530 86.920 99.620 91.430 ;
        RECT 100.890 91.240 101.300 91.320 ;
        RECT 90.530 77.570 94.550 86.920 ;
        RECT 99.900 86.060 100.140 91.050 ;
        RECT 100.290 91.010 101.300 91.240 ;
        RECT 100.890 90.940 101.300 91.010 ;
        RECT 100.300 89.950 100.710 90.020 ;
        RECT 100.290 89.720 101.290 89.950 ;
        RECT 100.300 89.640 100.710 89.720 ;
        RECT 100.890 88.660 101.300 88.730 ;
        RECT 100.290 88.430 101.300 88.660 ;
        RECT 100.890 88.350 101.300 88.430 ;
        RECT 100.290 87.370 100.700 87.450 ;
        RECT 100.290 87.140 101.290 87.370 ;
        RECT 100.290 87.070 100.700 87.140 ;
        RECT 101.440 86.060 101.680 91.050 ;
        RECT 113.010 87.220 113.280 93.040 ;
        RECT 114.970 91.750 115.630 91.840 ;
        RECT 113.475 91.520 115.630 91.750 ;
        RECT 114.970 91.440 115.630 91.520 ;
        RECT 113.480 91.110 114.140 91.200 ;
        RECT 113.475 90.880 115.615 91.110 ;
        RECT 113.480 90.800 114.140 90.880 ;
        RECT 114.970 90.470 115.630 90.560 ;
        RECT 113.475 90.240 115.630 90.470 ;
        RECT 114.970 90.160 115.630 90.240 ;
        RECT 113.480 89.830 114.140 89.910 ;
        RECT 113.475 89.600 115.615 89.830 ;
        RECT 113.480 89.510 114.140 89.600 ;
        RECT 114.970 89.190 115.630 89.280 ;
        RECT 113.475 88.960 115.630 89.190 ;
        RECT 114.970 88.880 115.630 88.960 ;
        RECT 113.470 88.550 114.130 88.640 ;
        RECT 113.470 88.320 115.615 88.550 ;
        RECT 113.470 88.240 114.130 88.320 ;
        RECT 114.970 87.910 115.630 88.000 ;
        RECT 113.475 87.680 115.630 87.910 ;
        RECT 114.970 87.600 115.630 87.680 ;
        RECT 113.480 87.270 114.140 87.360 ;
        RECT 113.475 87.040 115.615 87.270 ;
        RECT 115.800 87.220 116.070 93.040 ;
        RECT 118.930 91.960 120.090 100.150 ;
        RECT 116.330 90.800 120.090 91.960 ;
        RECT 113.480 86.960 114.140 87.040 ;
        RECT 116.330 86.800 117.780 90.800 ;
        RECT 99.900 85.970 101.680 86.060 ;
        RECT 103.825 85.970 104.555 86.000 ;
        RECT 99.900 85.240 104.555 85.970 ;
        RECT 123.350 85.350 123.580 116.340 ;
        RECT 125.190 114.970 125.790 115.050 ;
        RECT 123.785 114.740 125.790 114.970 ;
        RECT 125.190 114.660 125.790 114.740 ;
        RECT 123.790 111.680 124.390 111.760 ;
        RECT 123.785 111.450 125.785 111.680 ;
        RECT 123.790 111.370 124.390 111.450 ;
        RECT 125.190 108.390 125.790 108.470 ;
        RECT 123.785 108.160 125.790 108.390 ;
        RECT 125.190 108.080 125.790 108.160 ;
        RECT 123.790 105.100 124.390 105.190 ;
        RECT 123.785 104.870 125.785 105.100 ;
        RECT 123.790 104.800 124.390 104.870 ;
        RECT 125.190 101.810 125.790 101.900 ;
        RECT 123.785 101.580 125.790 101.810 ;
        RECT 125.190 101.510 125.790 101.580 ;
        RECT 123.790 98.520 124.390 98.600 ;
        RECT 123.785 98.290 125.785 98.520 ;
        RECT 123.790 98.210 124.390 98.290 ;
        RECT 125.190 95.230 125.790 95.310 ;
        RECT 123.785 95.000 125.790 95.230 ;
        RECT 125.190 94.920 125.790 95.000 ;
        RECT 123.790 91.940 124.390 92.020 ;
        RECT 123.785 91.710 125.785 91.940 ;
        RECT 123.790 91.630 124.390 91.710 ;
        RECT 125.190 88.650 125.790 88.740 ;
        RECT 123.785 88.420 125.790 88.650 ;
        RECT 125.190 88.350 125.790 88.420 ;
        RECT 123.790 85.360 124.390 85.440 ;
        RECT 99.900 85.200 101.680 85.240 ;
        RECT 103.825 85.210 104.555 85.240 ;
        RECT 123.785 85.130 125.785 85.360 ;
        RECT 125.990 85.350 126.220 116.340 ;
        RECT 128.600 115.190 132.620 120.240 ;
        RECT 123.790 85.050 124.390 85.130 ;
        RECT 126.500 84.900 132.620 115.190 ;
        RECT 96.720 82.935 98.295 82.965 ;
        RECT 100.430 82.935 110.130 82.940 ;
        RECT 96.720 81.400 110.130 82.935 ;
        RECT 128.600 82.160 132.620 84.900 ;
        RECT 125.120 81.460 132.620 82.160 ;
        RECT 96.720 81.360 102.285 81.400 ;
        RECT 96.720 81.330 98.295 81.360 ;
        RECT 97.975 77.570 98.705 79.795 ;
        RECT 128.600 79.695 132.620 81.460 ;
        RECT 126.025 79.005 132.620 79.695 ;
        RECT 99.930 78.370 106.195 78.880 ;
        RECT 90.530 72.870 99.640 77.570 ;
        RECT 99.930 73.390 100.170 78.370 ;
        RECT 100.320 77.270 100.690 77.350 ;
        RECT 100.320 77.040 101.320 77.270 ;
        RECT 100.320 76.970 100.690 77.040 ;
        RECT 100.950 75.980 101.320 76.060 ;
        RECT 100.320 75.750 101.320 75.980 ;
        RECT 100.950 75.680 101.320 75.750 ;
        RECT 100.310 74.690 100.680 74.770 ;
        RECT 100.310 74.460 101.320 74.690 ;
        RECT 100.310 74.390 100.680 74.460 ;
        RECT 100.950 73.400 101.320 73.480 ;
        RECT 100.320 73.170 101.320 73.400 ;
        RECT 101.460 73.390 101.730 78.370 ;
        RECT 100.950 73.100 101.320 73.170 ;
        RECT 90.530 69.585 94.550 72.870 ;
        RECT 112.720 71.310 113.890 78.980 ;
        RECT 115.160 78.720 115.560 78.810 ;
        RECT 114.560 78.490 115.560 78.720 ;
        RECT 90.530 69.330 110.805 69.585 ;
        RECT 112.720 69.330 113.620 71.310 ;
        RECT 114.160 70.640 114.410 78.480 ;
        RECT 115.160 78.410 115.560 78.490 ;
        RECT 114.550 76.430 114.950 76.520 ;
        RECT 114.550 76.200 115.560 76.430 ;
        RECT 114.550 76.120 114.950 76.200 ;
        RECT 115.170 74.140 115.570 74.230 ;
        RECT 114.560 73.910 115.570 74.140 ;
        RECT 115.170 73.830 115.570 73.910 ;
        RECT 114.550 71.850 114.950 71.940 ;
        RECT 114.550 71.620 115.560 71.850 ;
        RECT 114.550 71.540 114.950 71.620 ;
        RECT 115.710 70.640 115.960 78.480 ;
        RECT 128.600 78.140 132.620 79.005 ;
        RECT 124.600 77.890 125.110 77.970 ;
        RECT 123.435 77.660 125.110 77.890 ;
        RECT 120.895 75.415 121.945 76.405 ;
        RECT 120.925 71.635 121.915 75.415 ;
        RECT 122.980 74.460 123.260 77.660 ;
        RECT 124.600 77.580 125.110 77.660 ;
        RECT 123.450 77.250 123.960 77.330 ;
        RECT 123.435 77.020 125.105 77.250 ;
        RECT 123.450 76.940 123.960 77.020 ;
        RECT 124.600 76.610 125.110 76.690 ;
        RECT 123.435 76.380 125.110 76.610 ;
        RECT 124.600 76.300 125.110 76.380 ;
        RECT 123.450 75.970 123.960 76.050 ;
        RECT 123.435 75.740 125.105 75.970 ;
        RECT 123.450 75.660 123.960 75.740 ;
        RECT 125.290 74.460 125.570 77.660 ;
        RECT 125.800 75.460 132.620 78.140 ;
        RECT 122.980 74.180 125.570 74.460 ;
        RECT 123.030 72.800 123.310 74.180 ;
        RECT 120.925 70.645 125.685 71.635 ;
        RECT 114.160 70.050 115.960 70.640 ;
        RECT 90.530 68.430 113.620 69.330 ;
        RECT 115.160 69.950 115.960 70.050 ;
        RECT 122.780 70.590 125.680 70.645 ;
        RECT 115.160 68.930 119.490 69.950 ;
        RECT 90.530 68.175 110.805 68.430 ;
        RECT 90.530 45.450 94.550 68.175 ;
        RECT 111.570 66.120 112.310 66.800 ;
        RECT 101.800 64.120 103.010 64.130 ;
        RECT 104.040 64.120 104.725 66.050 ;
        RECT 105.900 65.280 111.265 65.290 ;
        RECT 111.600 65.280 112.280 66.120 ;
        RECT 105.640 64.860 113.930 65.280 ;
        RECT 101.800 62.890 105.450 64.120 ;
        RECT 105.640 63.290 105.930 64.860 ;
        RECT 106.090 63.850 106.500 63.940 ;
        RECT 106.090 63.620 107.090 63.850 ;
        RECT 106.090 63.570 106.500 63.620 ;
        RECT 106.680 63.410 107.090 63.470 ;
        RECT 106.090 63.180 107.090 63.410 ;
        RECT 107.240 63.290 107.530 64.860 ;
        RECT 110.980 63.240 111.270 64.860 ;
        RECT 112.850 63.900 113.470 63.980 ;
        RECT 111.465 63.670 113.470 63.900 ;
        RECT 112.850 63.600 113.470 63.670 ;
        RECT 111.480 63.260 112.100 63.340 ;
        RECT 106.680 63.100 107.090 63.180 ;
        RECT 111.465 63.030 113.465 63.260 ;
        RECT 113.640 63.240 113.930 64.860 ;
        RECT 114.825 64.180 115.720 66.165 ;
        RECT 111.480 62.960 112.100 63.030 ;
        RECT 101.800 59.440 104.580 62.890 ;
        RECT 114.150 62.770 117.250 64.180 ;
        RECT 109.000 61.240 109.685 62.415 ;
        RECT 105.900 61.230 113.940 61.240 ;
        RECT 105.670 60.800 113.940 61.230 ;
        RECT 105.670 60.780 111.270 60.800 ;
        RECT 101.800 57.730 105.430 59.440 ;
        RECT 105.670 58.620 105.950 60.780 ;
        RECT 107.120 59.170 107.550 59.250 ;
        RECT 106.090 58.940 107.590 59.170 ;
        RECT 107.120 58.850 107.550 58.940 ;
        RECT 106.140 58.690 106.570 58.770 ;
        RECT 106.090 58.460 107.590 58.690 ;
        RECT 106.140 58.370 106.570 58.460 ;
        RECT 107.120 58.210 107.550 58.300 ;
        RECT 106.090 57.980 107.590 58.210 ;
        RECT 107.730 58.140 108.020 60.780 ;
        RECT 107.120 57.900 107.550 57.980 ;
        RECT 110.980 57.850 111.260 60.780 ;
        RECT 112.900 59.760 113.460 59.850 ;
        RECT 111.465 59.530 113.465 59.760 ;
        RECT 112.900 59.450 113.460 59.530 ;
        RECT 111.480 59.120 112.040 59.200 ;
        RECT 111.465 58.890 113.465 59.120 ;
        RECT 111.480 58.800 112.040 58.890 ;
        RECT 112.900 58.480 113.460 58.570 ;
        RECT 111.465 58.250 113.465 58.480 ;
        RECT 112.900 58.170 113.460 58.250 ;
        RECT 111.480 57.840 112.040 57.920 ;
        RECT 113.650 57.850 113.930 60.800 ;
        RECT 115.330 60.030 117.250 62.770 ;
        RECT 101.800 52.600 103.010 57.730 ;
        RECT 111.465 57.610 113.465 57.840 ;
        RECT 111.480 57.520 112.040 57.610 ;
        RECT 114.140 57.340 117.250 60.030 ;
        RECT 104.030 55.540 106.420 56.220 ;
        RECT 108.925 55.540 109.800 57.040 ;
        RECT 104.030 55.520 111.385 55.540 ;
        RECT 104.030 54.850 114.920 55.520 ;
        RECT 104.030 54.830 111.385 54.850 ;
        RECT 104.030 54.675 106.420 54.830 ;
        RECT 101.800 50.410 103.990 52.600 ;
        RECT 104.230 50.840 104.500 54.675 ;
        RECT 104.710 52.340 105.220 52.440 ;
        RECT 104.650 52.110 107.650 52.340 ;
        RECT 104.710 52.010 105.220 52.110 ;
        RECT 107.090 51.860 107.600 51.960 ;
        RECT 104.650 51.630 107.650 51.860 ;
        RECT 107.090 51.530 107.600 51.630 ;
        RECT 104.720 51.380 105.230 51.480 ;
        RECT 104.650 51.150 107.650 51.380 ;
        RECT 107.800 51.320 108.070 54.830 ;
        RECT 104.720 51.050 105.230 51.150 ;
        RECT 107.090 50.900 107.600 51.000 ;
        RECT 104.650 50.670 107.650 50.900 ;
        RECT 107.090 50.570 107.600 50.670 ;
        RECT 101.800 45.450 103.460 50.410 ;
        RECT 110.980 49.680 111.260 54.830 ;
        RECT 113.860 53.540 114.460 53.620 ;
        RECT 111.465 53.310 114.465 53.540 ;
        RECT 113.860 53.220 114.460 53.310 ;
        RECT 111.500 52.900 112.100 52.980 ;
        RECT 111.465 52.670 114.465 52.900 ;
        RECT 111.500 52.580 112.100 52.670 ;
        RECT 113.860 52.260 114.460 52.350 ;
        RECT 111.465 52.030 114.465 52.260 ;
        RECT 113.860 51.950 114.460 52.030 ;
        RECT 111.500 51.620 112.100 51.710 ;
        RECT 111.465 51.390 114.465 51.620 ;
        RECT 111.500 51.310 112.100 51.390 ;
        RECT 113.860 50.980 114.460 51.060 ;
        RECT 111.465 50.750 114.465 50.980 ;
        RECT 113.860 50.660 114.460 50.750 ;
        RECT 111.500 50.340 112.100 50.430 ;
        RECT 111.465 50.110 114.465 50.340 ;
        RECT 111.500 50.030 112.100 50.110 ;
        RECT 113.860 49.700 114.460 49.790 ;
        RECT 111.465 49.470 114.465 49.700 ;
        RECT 114.640 49.680 114.920 54.850 ;
        RECT 116.100 53.740 117.250 57.340 ;
        RECT 113.860 49.390 114.460 49.470 ;
        RECT 115.170 49.220 117.250 53.740 ;
        RECT 118.470 52.550 119.490 68.930 ;
        RECT 90.530 43.790 103.460 45.450 ;
        RECT 108.480 45.155 109.560 47.520 ;
        RECT 115.440 45.275 117.250 49.220 ;
        RECT 118.150 48.725 119.615 52.550 ;
        RECT 122.780 49.580 123.040 70.590 ;
        RECT 123.250 69.330 123.820 69.430 ;
        RECT 123.235 69.100 125.235 69.330 ;
        RECT 123.250 69.010 123.820 69.100 ;
        RECT 124.670 66.040 125.240 66.140 ;
        RECT 123.235 65.810 125.240 66.040 ;
        RECT 124.670 65.720 125.240 65.810 ;
        RECT 123.250 62.750 123.820 62.860 ;
        RECT 123.235 62.520 125.235 62.750 ;
        RECT 123.250 62.440 123.820 62.520 ;
        RECT 124.680 59.460 125.250 59.560 ;
        RECT 123.235 59.230 125.250 59.460 ;
        RECT 124.680 59.140 125.250 59.230 ;
        RECT 123.250 56.170 123.820 56.270 ;
        RECT 123.235 55.940 125.235 56.170 ;
        RECT 123.250 55.850 123.820 55.940 ;
        RECT 124.680 52.880 125.250 52.980 ;
        RECT 123.235 52.650 125.250 52.880 ;
        RECT 124.680 52.560 125.250 52.650 ;
        RECT 123.250 49.590 123.820 49.680 ;
        RECT 123.235 49.360 125.235 49.590 ;
        RECT 125.420 49.580 125.680 70.590 ;
        RECT 128.600 69.590 132.620 75.460 ;
        RECT 123.250 49.260 123.820 49.360 ;
        RECT 125.960 49.060 132.620 69.590 ;
        RECT 118.120 47.260 119.645 48.725 ;
        RECT 128.600 47.555 132.620 49.060 ;
        RECT 124.555 46.740 132.620 47.555 ;
        RECT 128.600 45.275 132.620 46.740 ;
        RECT 90.530 42.990 94.550 43.790 ;
        RECT 108.045 38.585 109.660 45.155 ;
        RECT 115.440 43.465 132.620 45.275 ;
        RECT 128.600 42.990 132.620 43.465 ;
        RECT 108.015 36.970 109.690 38.585 ;
      LAYER via ;
        RECT 129.155 159.540 131.840 162.225 ;
        RECT 87.860 151.120 89.820 153.080 ;
        RECT 118.920 146.110 120.300 147.490 ;
        RECT 103.490 131.920 104.050 132.480 ;
        RECT 108.830 136.880 109.320 137.170 ;
        RECT 106.390 136.420 106.880 136.710 ;
        RECT 108.830 135.940 109.320 136.230 ;
        RECT 106.390 135.460 106.880 135.750 ;
        RECT 108.830 134.980 109.320 135.270 ;
        RECT 106.390 134.500 106.880 134.790 ;
        RECT 108.830 134.020 109.320 134.310 ;
        RECT 106.390 133.540 106.880 133.830 ;
        RECT 108.015 131.970 108.585 132.540 ;
        RECT 111.750 133.410 113.315 134.975 ;
        RECT 115.570 136.840 116.050 137.120 ;
        RECT 117.970 136.270 118.450 136.550 ;
        RECT 115.550 135.620 116.030 135.900 ;
        RECT 117.970 134.980 118.450 135.260 ;
        RECT 115.550 134.350 116.030 134.630 ;
        RECT 117.970 133.710 118.450 133.990 ;
        RECT 115.550 133.060 116.030 133.340 ;
        RECT 117.970 132.430 118.450 132.710 ;
        RECT 115.520 130.710 116.100 131.290 ;
        RECT 125.630 127.755 126.220 128.345 ;
        RECT 100.540 121.710 101.170 122.030 ;
        RECT 97.310 118.440 97.940 118.760 ;
        RECT 100.540 115.130 101.170 115.450 ;
        RECT 97.310 111.830 97.940 112.150 ;
        RECT 97.260 109.770 98.010 110.520 ;
        RECT 100.540 106.080 101.250 106.450 ;
        RECT 97.360 102.790 98.070 103.160 ;
        RECT 100.540 99.510 101.250 99.880 ;
        RECT 97.360 96.220 98.070 96.590 ;
        RECT 109.150 118.080 109.560 118.370 ;
        RECT 108.170 117.090 108.580 117.380 ;
        RECT 109.150 116.100 109.560 116.390 ;
        RECT 108.170 115.110 108.580 115.400 ;
        RECT 109.150 114.120 109.560 114.410 ;
        RECT 108.170 113.130 108.580 113.420 ;
        RECT 109.150 112.140 109.560 112.430 ;
        RECT 108.170 111.160 108.580 111.450 ;
        RECT 109.150 110.160 109.560 110.450 ;
        RECT 108.170 109.180 108.580 109.470 ;
        RECT 109.150 108.180 109.560 108.470 ;
        RECT 108.170 107.190 108.580 107.480 ;
        RECT 109.150 106.200 109.560 106.490 ;
        RECT 108.170 105.220 108.580 105.510 ;
        RECT 109.150 104.220 109.560 104.510 ;
        RECT 108.170 103.230 108.580 103.520 ;
        RECT 109.150 102.240 109.560 102.530 ;
        RECT 108.170 101.250 108.580 101.540 ;
        RECT 109.150 100.260 109.560 100.550 ;
        RECT 116.940 118.080 117.470 118.370 ;
        RECT 115.980 117.090 116.510 117.380 ;
        RECT 116.940 116.100 117.470 116.390 ;
        RECT 115.980 115.120 116.510 115.410 ;
        RECT 116.940 114.120 117.470 114.410 ;
        RECT 115.980 113.140 116.510 113.430 ;
        RECT 116.940 112.150 117.470 112.440 ;
        RECT 115.980 111.150 116.510 111.440 ;
        RECT 116.940 110.170 117.470 110.460 ;
        RECT 115.980 109.170 116.510 109.460 ;
        RECT 116.940 108.180 117.470 108.470 ;
        RECT 115.980 107.200 116.510 107.490 ;
        RECT 116.940 106.200 117.470 106.490 ;
        RECT 115.980 105.220 116.510 105.510 ;
        RECT 116.940 104.230 117.470 104.520 ;
        RECT 115.980 103.240 116.510 103.530 ;
        RECT 116.940 102.240 117.470 102.530 ;
        RECT 115.980 101.260 116.510 101.550 ;
        RECT 116.940 100.260 117.470 100.550 ;
        RECT 125.630 117.365 126.220 117.955 ;
        RECT 106.435 95.785 107.125 96.475 ;
        RECT 97.320 93.790 98.120 94.590 ;
        RECT 113.010 94.435 113.680 95.105 ;
        RECT 100.340 92.320 100.700 92.680 ;
        RECT 100.890 90.990 101.300 91.270 ;
        RECT 100.300 89.690 100.710 89.970 ;
        RECT 100.890 88.400 101.300 88.680 ;
        RECT 100.290 87.120 100.700 87.400 ;
        RECT 114.970 91.490 115.630 91.790 ;
        RECT 113.480 90.850 114.140 91.150 ;
        RECT 114.970 90.210 115.630 90.510 ;
        RECT 113.480 89.560 114.140 89.860 ;
        RECT 114.970 88.930 115.630 89.230 ;
        RECT 113.470 88.290 114.130 88.590 ;
        RECT 114.970 87.650 115.630 87.950 ;
        RECT 113.480 87.010 114.140 87.310 ;
        RECT 100.950 85.515 101.340 85.905 ;
        RECT 103.825 85.240 104.555 85.970 ;
        RECT 125.190 114.710 125.790 115.000 ;
        RECT 123.790 111.420 124.390 111.710 ;
        RECT 125.190 108.130 125.790 108.420 ;
        RECT 123.790 104.850 124.390 105.140 ;
        RECT 125.190 101.560 125.790 101.850 ;
        RECT 123.790 98.260 124.390 98.550 ;
        RECT 125.190 94.970 125.790 95.260 ;
        RECT 123.790 91.680 124.390 91.970 ;
        RECT 125.190 88.400 125.790 88.690 ;
        RECT 123.790 85.100 124.390 85.390 ;
        RECT 108.560 81.400 110.100 82.940 ;
        RECT 125.150 81.460 125.850 82.160 ;
        RECT 97.975 79.035 98.705 79.765 ;
        RECT 126.080 79.060 126.660 79.640 ;
        RECT 105.655 78.370 106.165 78.880 ;
        RECT 100.320 77.020 100.690 77.300 ;
        RECT 100.950 75.730 101.320 76.010 ;
        RECT 100.310 74.440 100.680 74.720 ;
        RECT 100.950 73.150 101.320 73.430 ;
        RECT 115.160 78.460 115.560 78.760 ;
        RECT 114.550 76.170 114.950 76.470 ;
        RECT 115.170 73.880 115.570 74.180 ;
        RECT 114.550 71.590 114.950 71.890 ;
        RECT 120.925 75.415 121.915 76.405 ;
        RECT 124.600 77.630 125.110 77.920 ;
        RECT 123.450 76.990 123.960 77.280 ;
        RECT 124.600 76.350 125.110 76.640 ;
        RECT 123.450 75.710 123.960 76.000 ;
        RECT 123.030 72.830 123.310 73.110 ;
        RECT 111.600 66.120 112.280 66.800 ;
        RECT 104.125 65.455 104.635 65.965 ;
        RECT 114.905 65.355 115.635 66.085 ;
        RECT 106.680 63.150 107.090 63.420 ;
        RECT 112.850 63.650 113.470 63.930 ;
        RECT 111.480 63.010 112.100 63.290 ;
        RECT 109.075 61.810 109.605 62.340 ;
        RECT 103.430 59.980 103.950 60.500 ;
        RECT 115.735 60.925 116.385 61.575 ;
        RECT 107.120 58.900 107.550 59.200 ;
        RECT 106.140 58.420 106.570 58.720 ;
        RECT 107.120 57.950 107.550 58.250 ;
        RECT 112.900 59.500 113.460 59.800 ;
        RECT 111.480 58.850 112.040 59.150 ;
        RECT 112.900 58.220 113.460 58.520 ;
        RECT 111.480 57.570 112.040 57.870 ;
        RECT 109.035 56.280 109.685 56.930 ;
        RECT 104.235 54.885 105.365 56.015 ;
        RECT 104.710 52.060 105.220 52.390 ;
        RECT 107.090 51.580 107.600 51.910 ;
        RECT 104.720 51.100 105.230 51.430 ;
        RECT 107.090 50.620 107.600 50.950 ;
        RECT 113.860 53.270 114.460 53.570 ;
        RECT 111.500 52.630 112.100 52.930 ;
        RECT 113.860 52.000 114.460 52.300 ;
        RECT 111.500 51.360 112.100 51.660 ;
        RECT 113.860 50.710 114.460 51.010 ;
        RECT 111.500 50.080 112.100 50.380 ;
        RECT 113.860 49.440 114.460 49.740 ;
        RECT 102.445 48.580 103.075 49.210 ;
        RECT 123.250 69.060 123.820 69.380 ;
        RECT 124.670 65.770 125.240 66.090 ;
        RECT 123.250 62.490 123.820 62.810 ;
        RECT 124.680 59.190 125.250 59.510 ;
        RECT 123.250 55.900 123.820 56.220 ;
        RECT 124.680 52.610 125.250 52.930 ;
        RECT 123.250 49.310 123.820 49.630 ;
        RECT 115.855 47.600 116.625 48.370 ;
        RECT 108.705 46.665 109.335 47.295 ;
        RECT 118.150 47.260 119.615 48.725 ;
        RECT 124.640 46.830 125.280 47.470 ;
        RECT 108.045 36.970 109.660 38.585 ;
      LAYER met2 ;
        RECT 129.155 162.225 131.840 162.255 ;
        RECT 79.225 161.760 80.910 161.770 ;
        RECT 87.495 161.760 131.840 162.225 ;
        RECT 79.190 160.005 131.840 161.760 ;
        RECT 79.225 159.995 80.910 160.005 ;
        RECT 87.495 159.540 131.840 160.005 ;
        RECT 129.155 159.510 131.840 159.540 ;
        RECT 75.895 152.850 77.345 152.870 ;
        RECT 83.160 152.850 89.850 153.080 ;
        RECT 75.870 151.350 89.850 152.850 ;
        RECT 75.895 151.330 77.345 151.350 ;
        RECT 83.160 151.120 89.850 151.350 ;
        RECT 121.325 147.490 122.655 147.510 ;
        RECT 118.890 146.110 122.680 147.490 ;
        RECT 121.325 146.090 122.655 146.110 ;
        RECT 108.780 136.880 109.370 137.170 ;
        RECT 106.340 136.420 106.930 136.710 ;
        RECT 106.370 135.750 106.930 136.420 ;
        RECT 108.800 136.230 109.370 136.880 ;
        RECT 108.780 135.940 109.370 136.230 ;
        RECT 106.340 135.460 106.930 135.750 ;
        RECT 106.370 134.790 106.930 135.460 ;
        RECT 108.800 135.270 109.370 135.940 ;
        RECT 115.520 135.900 116.100 137.130 ;
        RECT 117.940 136.550 118.480 136.610 ;
        RECT 117.920 136.270 118.500 136.550 ;
        RECT 115.500 135.620 116.100 135.900 ;
        RECT 108.780 134.980 109.370 135.270 ;
        RECT 106.340 134.500 106.930 134.790 ;
        RECT 106.370 133.830 106.930 134.500 ;
        RECT 108.800 134.310 109.370 134.980 ;
        RECT 108.780 134.020 109.370 134.310 ;
        RECT 106.340 133.540 106.930 133.830 ;
        RECT 103.490 132.480 104.050 132.510 ;
        RECT 106.370 132.480 106.930 133.540 ;
        RECT 108.800 132.540 109.370 134.020 ;
        RECT 111.720 133.410 113.345 134.975 ;
        RECT 115.520 134.630 116.100 135.620 ;
        RECT 117.940 135.260 118.480 136.270 ;
        RECT 117.920 134.980 118.500 135.260 ;
        RECT 115.500 134.350 116.100 134.630 ;
        RECT 103.490 131.920 106.930 132.480 ;
        RECT 107.985 131.970 109.370 132.540 ;
        RECT 103.490 131.890 104.050 131.920 ;
        RECT 111.750 125.765 113.315 133.410 ;
        RECT 115.520 133.340 116.100 134.350 ;
        RECT 117.940 133.990 118.480 134.980 ;
        RECT 117.920 133.710 118.500 133.990 ;
        RECT 115.500 133.060 116.100 133.340 ;
        RECT 115.520 130.680 116.100 133.060 ;
        RECT 117.940 132.710 118.480 133.710 ;
        RECT 117.920 132.430 118.500 132.710 ;
        RECT 117.940 131.250 118.480 132.430 ;
        RECT 117.940 130.710 121.010 131.250 ;
        RECT 100.490 123.560 109.705 124.270 ;
        RECT 111.750 124.200 117.960 125.765 ;
        RECT 100.490 122.030 101.200 123.560 ;
        RECT 100.490 121.710 101.220 122.030 ;
        RECT 97.260 109.740 98.010 118.830 ;
        RECT 100.490 115.450 101.200 121.710 ;
        RECT 108.995 121.185 109.705 123.560 ;
        RECT 116.395 122.050 117.960 124.200 ;
        RECT 115.940 121.185 116.530 121.210 ;
        RECT 108.995 120.475 116.530 121.185 ;
        RECT 109.110 118.370 109.620 118.420 ;
        RECT 109.100 118.080 109.620 118.370 ;
        RECT 100.490 115.130 101.220 115.450 ;
        RECT 100.490 114.730 101.200 115.130 ;
        RECT 100.470 106.450 101.270 106.560 ;
        RECT 100.470 106.080 101.300 106.450 ;
        RECT 97.320 103.160 98.120 103.270 ;
        RECT 97.310 102.790 98.120 103.160 ;
        RECT 97.320 96.590 98.120 102.790 ;
        RECT 97.310 96.220 98.120 96.590 ;
        RECT 97.320 93.760 98.120 96.220 ;
        RECT 100.470 99.880 101.270 106.080 ;
        RECT 100.470 99.510 101.300 99.880 ;
        RECT 100.470 94.780 101.270 99.510 ;
        RECT 108.060 96.640 108.720 117.580 ;
        RECT 109.110 116.390 109.620 118.080 ;
        RECT 109.100 116.100 109.620 116.390 ;
        RECT 109.110 114.410 109.620 116.100 ;
        RECT 109.100 114.120 109.620 114.410 ;
        RECT 109.110 112.430 109.620 114.120 ;
        RECT 109.100 112.140 109.620 112.430 ;
        RECT 109.110 110.450 109.620 112.140 ;
        RECT 109.100 110.160 109.620 110.450 ;
        RECT 109.110 108.470 109.620 110.160 ;
        RECT 109.100 108.180 109.620 108.470 ;
        RECT 109.110 106.490 109.620 108.180 ;
        RECT 109.100 106.200 109.620 106.490 ;
        RECT 109.110 104.510 109.620 106.200 ;
        RECT 109.100 104.220 109.620 104.510 ;
        RECT 109.110 102.530 109.620 104.220 ;
        RECT 109.100 102.240 109.620 102.530 ;
        RECT 109.110 100.550 109.620 102.240 ;
        RECT 109.100 100.260 109.620 100.550 ;
        RECT 108.060 96.475 108.750 96.640 ;
        RECT 106.405 95.785 108.750 96.475 ;
        RECT 108.060 95.580 108.750 95.785 ;
        RECT 108.060 94.780 108.720 95.580 ;
        RECT 100.470 93.980 108.790 94.780 ;
        RECT 109.110 93.575 109.620 100.260 ;
        RECT 113.010 95.105 113.680 120.475 ;
        RECT 115.940 117.380 116.530 120.475 ;
        RECT 116.840 118.370 117.510 122.050 ;
        RECT 120.925 118.995 121.915 119.195 ;
        RECT 125.630 118.995 126.220 128.375 ;
        RECT 120.925 118.405 126.220 118.995 ;
        RECT 116.840 118.080 117.520 118.370 ;
        RECT 115.930 117.090 116.560 117.380 ;
        RECT 115.940 115.410 116.530 117.090 ;
        RECT 116.840 116.390 117.510 118.080 ;
        RECT 116.840 116.100 117.520 116.390 ;
        RECT 115.930 115.120 116.560 115.410 ;
        RECT 115.940 113.430 116.530 115.120 ;
        RECT 116.840 114.410 117.510 116.100 ;
        RECT 116.840 114.120 117.520 114.410 ;
        RECT 115.930 113.140 116.560 113.430 ;
        RECT 115.940 111.440 116.530 113.140 ;
        RECT 116.840 112.440 117.510 114.120 ;
        RECT 116.840 112.150 117.520 112.440 ;
        RECT 115.930 111.150 116.560 111.440 ;
        RECT 115.940 109.460 116.530 111.150 ;
        RECT 116.840 110.460 117.510 112.150 ;
        RECT 116.840 110.170 117.520 110.460 ;
        RECT 115.930 109.170 116.560 109.460 ;
        RECT 115.940 107.490 116.530 109.170 ;
        RECT 116.840 108.470 117.510 110.170 ;
        RECT 116.840 108.180 117.520 108.470 ;
        RECT 115.930 107.200 116.560 107.490 ;
        RECT 115.940 105.510 116.530 107.200 ;
        RECT 116.840 106.490 117.510 108.180 ;
        RECT 116.840 106.200 117.520 106.490 ;
        RECT 115.930 105.220 116.560 105.510 ;
        RECT 115.940 103.530 116.530 105.220 ;
        RECT 116.840 104.520 117.510 106.200 ;
        RECT 116.840 104.230 117.520 104.520 ;
        RECT 115.930 103.240 116.560 103.530 ;
        RECT 115.940 101.550 116.530 103.240 ;
        RECT 116.840 102.530 117.510 104.230 ;
        RECT 116.840 102.240 117.520 102.530 ;
        RECT 115.930 101.260 116.560 101.550 ;
        RECT 115.940 101.140 116.530 101.260 ;
        RECT 116.840 100.550 117.510 102.240 ;
        RECT 116.840 100.260 117.520 100.550 ;
        RECT 116.840 100.225 117.510 100.260 ;
        RECT 112.980 94.435 113.710 95.105 ;
        RECT 109.110 93.065 119.405 93.575 ;
        RECT 100.310 92.320 100.730 92.680 ;
        RECT 100.340 89.970 100.700 92.320 ;
        RECT 100.840 90.990 101.350 91.270 ;
        RECT 113.490 91.150 114.220 91.200 ;
        RECT 100.250 89.690 100.760 89.970 ;
        RECT 100.340 87.400 100.700 89.690 ;
        RECT 100.950 88.680 101.340 90.990 ;
        RECT 113.430 90.850 114.220 91.150 ;
        RECT 113.490 89.860 114.220 90.850 ;
        RECT 113.430 89.560 114.220 89.860 ;
        RECT 100.840 88.400 101.350 88.680 ;
        RECT 113.490 88.590 114.220 89.560 ;
        RECT 100.240 87.120 100.750 87.400 ;
        RECT 100.340 87.110 100.700 87.120 ;
        RECT 100.950 85.485 101.340 88.400 ;
        RECT 113.420 88.290 114.220 88.590 ;
        RECT 113.490 87.310 114.220 88.290 ;
        RECT 114.910 87.500 115.680 93.065 ;
        RECT 113.430 87.010 114.220 87.310 ;
        RECT 113.490 85.970 114.220 87.010 ;
        RECT 103.795 85.240 114.220 85.970 ;
        RECT 75.235 81.360 98.325 82.935 ;
        RECT 75.235 67.550 76.810 81.360 ;
        RECT 97.945 79.630 99.415 79.765 ;
        RECT 97.945 79.170 100.730 79.630 ;
        RECT 97.945 79.035 99.415 79.170 ;
        RECT 100.270 77.300 100.730 79.170 ;
        RECT 105.510 78.220 106.315 85.240 ;
        RECT 118.895 84.805 119.405 93.065 ;
        RECT 120.925 86.720 121.915 118.405 ;
        RECT 125.630 117.955 126.220 118.405 ;
        RECT 125.600 117.365 126.250 117.955 ;
        RECT 125.150 115.000 125.850 115.060 ;
        RECT 125.140 114.710 125.850 115.000 ;
        RECT 123.750 111.710 124.450 111.810 ;
        RECT 123.740 111.420 124.450 111.710 ;
        RECT 123.750 105.140 124.450 111.420 ;
        RECT 125.150 108.420 125.850 114.710 ;
        RECT 125.140 108.130 125.850 108.420 ;
        RECT 123.740 104.850 124.450 105.140 ;
        RECT 123.750 98.550 124.450 104.850 ;
        RECT 125.150 101.850 125.850 108.130 ;
        RECT 125.140 101.560 125.850 101.850 ;
        RECT 123.740 98.260 124.450 98.550 ;
        RECT 123.750 91.970 124.450 98.260 ;
        RECT 125.150 95.260 125.850 101.560 ;
        RECT 125.140 94.970 125.850 95.260 ;
        RECT 123.740 91.680 124.450 91.970 ;
        RECT 123.750 85.390 124.450 91.680 ;
        RECT 125.150 88.690 125.850 94.970 ;
        RECT 125.140 88.400 125.850 88.690 ;
        RECT 123.740 85.100 124.450 85.390 ;
        RECT 118.885 84.235 119.405 84.805 ;
        RECT 118.885 83.300 119.395 84.235 ;
        RECT 123.750 83.300 124.450 85.100 ;
        RECT 108.560 82.940 110.100 82.970 ;
        RECT 108.560 82.910 114.970 82.940 ;
        RECT 118.880 82.910 124.450 83.300 ;
        RECT 108.560 81.465 124.450 82.910 ;
        RECT 108.560 81.400 114.970 81.465 ;
        RECT 118.880 81.460 124.450 81.465 ;
        RECT 125.150 81.430 125.850 88.400 ;
        RECT 108.560 81.370 110.100 81.400 ;
        RECT 100.270 77.020 100.740 77.300 ;
        RECT 100.270 74.720 100.730 77.020 ;
        RECT 114.490 76.470 114.950 81.400 ;
        RECT 115.160 79.670 124.000 80.120 ;
        RECT 115.160 78.760 115.610 79.670 ;
        RECT 115.110 78.460 115.610 78.760 ;
        RECT 114.490 76.170 115.000 76.470 ;
        RECT 100.920 76.010 101.370 76.040 ;
        RECT 100.900 75.730 101.370 76.010 ;
        RECT 100.260 74.440 100.730 74.720 ;
        RECT 100.270 74.410 100.730 74.440 ;
        RECT 100.920 73.430 101.370 75.730 ;
        RECT 100.900 73.150 101.370 73.430 ;
        RECT 100.920 71.370 101.370 73.150 ;
        RECT 114.490 71.890 114.950 76.170 ;
        RECT 115.160 74.180 115.610 78.460 ;
        RECT 120.925 77.850 121.915 77.875 ;
        RECT 115.120 73.880 115.620 74.180 ;
        RECT 118.345 73.955 119.475 77.840 ;
        RECT 120.905 76.910 121.935 77.850 ;
        RECT 123.390 77.280 124.000 79.670 ;
        RECT 124.580 79.060 126.690 79.640 ;
        RECT 124.580 77.920 125.160 79.060 ;
        RECT 124.550 77.630 125.160 77.920 ;
        RECT 123.390 76.990 124.010 77.280 ;
        RECT 120.925 75.385 121.915 76.910 ;
        RECT 123.390 76.000 124.000 76.990 ;
        RECT 124.580 76.640 125.160 77.630 ;
        RECT 124.550 76.350 125.160 76.640 ;
        RECT 124.580 76.310 125.160 76.350 ;
        RECT 123.390 75.710 124.010 76.000 ;
        RECT 123.390 75.690 124.000 75.710 ;
        RECT 115.160 73.780 115.610 73.880 ;
        RECT 118.600 73.280 119.225 73.955 ;
        RECT 118.600 72.655 123.485 73.280 ;
        RECT 114.490 71.590 115.000 71.890 ;
        RECT 114.490 71.550 114.950 71.590 ;
        RECT 100.920 70.105 112.280 71.370 ;
        RECT 101.300 70.080 112.280 70.105 ;
        RECT 111.590 68.020 112.270 70.080 ;
        RECT 75.215 66.025 76.830 67.550 ;
        RECT 111.590 67.430 117.130 68.020 ;
        RECT 111.590 67.415 119.730 67.430 ;
        RECT 111.590 67.340 121.725 67.415 ;
        RECT 111.600 66.090 112.280 67.340 ;
        RECT 116.450 66.750 121.725 67.340 ;
        RECT 119.185 66.725 121.725 66.750 ;
        RECT 75.235 66.000 76.810 66.025 ;
        RECT 104.095 65.455 106.550 65.965 ;
        RECT 106.040 63.620 106.550 65.455 ;
        RECT 112.800 65.355 115.665 66.085 ;
        RECT 112.800 63.650 113.530 65.355 ;
        RECT 106.630 62.340 107.160 63.420 ;
        RECT 111.420 62.340 112.150 63.300 ;
        RECT 106.630 61.810 112.150 62.340 ;
        RECT 112.860 60.925 116.415 61.575 ;
        RECT 103.400 59.980 106.610 60.500 ;
        RECT 106.090 58.720 106.610 59.980 ;
        RECT 112.860 59.800 113.510 60.925 ;
        RECT 112.850 59.500 113.510 59.800 ;
        RECT 107.100 59.200 107.600 59.220 ;
        RECT 107.070 58.900 107.600 59.200 ;
        RECT 106.090 58.420 106.620 58.720 ;
        RECT 106.090 58.390 106.610 58.420 ;
        RECT 107.100 58.250 107.600 58.900 ;
        RECT 107.070 57.950 107.600 58.250 ;
        RECT 107.100 56.930 107.600 57.950 ;
        RECT 111.430 59.150 112.080 59.190 ;
        RECT 111.430 58.850 112.090 59.150 ;
        RECT 111.430 57.870 112.080 58.850 ;
        RECT 112.860 58.520 113.510 59.500 ;
        RECT 112.850 58.220 113.510 58.520 ;
        RECT 112.860 58.200 113.510 58.220 ;
        RECT 111.430 57.570 112.090 57.870 ;
        RECT 109.035 56.930 109.685 56.960 ;
        RECT 111.430 56.930 112.080 57.570 ;
        RECT 107.095 56.280 112.080 56.930 ;
        RECT 107.100 56.260 107.600 56.280 ;
        RECT 109.035 56.250 109.685 56.280 ;
        RECT 98.575 55.990 105.395 56.015 ;
        RECT 98.555 54.910 105.395 55.990 ;
        RECT 98.575 54.885 105.395 54.910 ;
        RECT 104.650 49.210 105.280 52.440 ;
        RECT 102.415 48.580 105.280 49.210 ;
        RECT 107.020 48.220 107.650 51.920 ;
        RECT 111.450 48.220 112.160 52.940 ;
        RECT 107.020 47.590 112.160 48.220 ;
        RECT 113.750 48.370 114.520 53.630 ;
        RECT 113.750 47.600 116.655 48.370 ;
        RECT 108.705 46.635 109.335 47.590 ;
        RECT 118.150 38.825 119.615 48.755 ;
        RECT 121.035 48.200 121.725 66.725 ;
        RECT 123.180 48.200 123.870 69.440 ;
        RECT 124.640 66.090 125.280 66.180 ;
        RECT 124.620 65.770 125.290 66.090 ;
        RECT 124.640 59.510 125.280 65.770 ;
        RECT 124.630 59.190 125.300 59.510 ;
        RECT 124.640 52.930 125.280 59.190 ;
        RECT 124.630 52.610 125.300 52.930 ;
        RECT 121.035 47.510 123.870 48.200 ;
        RECT 124.640 47.470 125.280 52.610 ;
        RECT 124.610 46.830 125.310 47.470 ;
        RECT 108.045 33.220 109.660 38.615 ;
        RECT 118.130 37.410 119.635 38.825 ;
        RECT 118.150 37.385 119.615 37.410 ;
        RECT 108.025 31.655 109.680 33.220 ;
        RECT 108.045 31.630 109.660 31.655 ;
      LAYER via2 ;
        RECT 79.225 160.040 80.910 161.725 ;
        RECT 75.895 151.375 77.345 152.825 ;
        RECT 121.325 146.135 122.655 147.465 ;
        RECT 120.925 86.765 121.915 87.755 ;
        RECT 118.345 76.665 119.475 77.795 ;
        RECT 120.950 76.910 121.890 77.850 ;
        RECT 75.260 66.025 76.785 67.550 ;
        RECT 98.600 54.910 99.680 55.990 ;
        RECT 118.175 37.410 119.590 38.825 ;
        RECT 108.070 31.655 109.635 33.220 ;
      LAYER met3 ;
        RECT 30.455 161.630 31.945 161.655 ;
        RECT 74.815 161.630 80.935 161.750 ;
        RECT 30.450 160.130 80.935 161.630 ;
        RECT 30.455 160.105 31.945 160.130 ;
        RECT 74.815 160.015 80.935 160.130 ;
        RECT 71.175 152.850 72.665 152.875 ;
        RECT 71.170 151.350 77.370 152.850 ;
        RECT 71.175 151.325 72.665 151.350 ;
        RECT 123.835 147.490 125.205 147.515 ;
        RECT 121.300 146.110 125.210 147.490 ;
        RECT 123.835 146.085 125.205 146.110 ;
        RECT 120.900 86.740 121.940 87.780 ;
        RECT 110.825 80.545 119.475 81.675 ;
        RECT 110.825 74.935 111.955 80.545 ;
        RECT 118.345 77.820 119.475 80.545 ;
        RECT 118.320 76.640 119.500 77.820 ;
        RECT 120.925 76.885 121.915 86.740 ;
        RECT 104.855 73.805 111.955 74.935 ;
        RECT 104.855 69.035 105.985 73.805 ;
        RECT 98.575 67.905 105.985 69.035 ;
        RECT 75.235 59.600 76.810 67.575 ;
        RECT 75.210 58.035 76.835 59.600 ;
        RECT 75.235 58.030 76.810 58.035 ;
        RECT 98.575 54.885 99.705 67.905 ;
        RECT 118.150 33.675 119.615 38.850 ;
        RECT 108.045 28.040 109.660 33.245 ;
        RECT 118.125 32.220 119.640 33.675 ;
        RECT 118.150 32.215 119.615 32.220 ;
        RECT 108.020 26.435 109.685 28.040 ;
        RECT 108.045 26.430 109.660 26.435 ;
      LAYER via3 ;
        RECT 30.455 160.135 31.945 161.625 ;
        RECT 71.175 151.355 72.665 152.845 ;
        RECT 123.835 146.115 125.205 147.485 ;
        RECT 75.240 58.035 76.805 59.600 ;
        RECT 118.155 32.220 119.610 33.675 ;
        RECT 108.050 26.435 109.655 28.040 ;
      LAYER met4 ;
        RECT 3.990 223.570 4.290 224.760 ;
        RECT 7.670 223.570 7.970 224.760 ;
        RECT 11.350 223.570 11.650 224.760 ;
        RECT 15.030 223.570 15.330 224.760 ;
        RECT 18.710 223.570 19.010 224.760 ;
        RECT 22.390 223.570 22.690 224.760 ;
        RECT 26.070 223.570 26.370 224.760 ;
        RECT 29.750 223.570 30.050 224.760 ;
        RECT 33.430 223.570 33.730 224.760 ;
        RECT 37.110 223.570 37.410 224.760 ;
        RECT 40.790 223.570 41.090 224.760 ;
        RECT 44.470 223.570 44.770 224.760 ;
        RECT 48.150 223.570 48.450 224.760 ;
        RECT 51.830 223.570 52.130 224.760 ;
        RECT 55.510 223.570 55.810 224.760 ;
        RECT 59.190 223.570 59.490 224.760 ;
        RECT 62.870 223.570 63.170 224.760 ;
        RECT 66.550 223.570 66.850 224.760 ;
        RECT 70.230 223.570 70.530 224.760 ;
        RECT 73.910 223.570 74.210 224.760 ;
        RECT 77.590 223.570 77.890 224.760 ;
        RECT 81.270 223.570 81.570 224.760 ;
        RECT 84.950 223.570 85.250 224.760 ;
        RECT 88.630 223.570 88.930 224.760 ;
        RECT 3.760 222.150 88.940 223.570 ;
        RECT 49.000 220.760 50.500 222.150 ;
        RECT 2.500 160.130 31.950 161.630 ;
        RECT 50.500 151.350 72.670 152.850 ;
        RECT 123.830 146.110 145.730 147.490 ;
        RECT 75.235 23.435 76.810 59.605 ;
        RECT 118.150 32.215 135.515 33.680 ;
        RECT 75.235 21.860 91.410 23.435 ;
        RECT 89.835 8.495 91.410 21.860 ;
        RECT 108.045 21.625 109.660 28.045 ;
        RECT 108.045 20.010 113.510 21.625 ;
        RECT 111.895 9.775 113.510 20.010 ;
        RECT 134.050 17.240 135.515 32.215 ;
        RECT 144.350 17.980 145.730 146.110 ;
        RECT 144.350 17.590 152.430 17.980 ;
        RECT 156.560 17.590 157.160 17.660 ;
        RECT 90.320 1.000 90.920 8.495 ;
        RECT 112.400 1.000 113.000 9.775 ;
        RECT 134.480 1.000 135.080 17.240 ;
        RECT 144.350 16.990 157.160 17.590 ;
        RECT 144.350 16.600 152.430 16.990 ;
        RECT 156.560 1.000 157.160 16.990 ;
  END
END tt_um_alfiero88_CurrentTrigger
END LIBRARY


magic
tech sky130A
magscale 1 2
timestamp 1717082428
<< viali >>
rect 246 9102 982 9142
rect 4660 8882 10668 8930
rect 12072 8746 12546 8796
rect 13786 8774 17822 8822
rect 126 6584 166 7364
rect 4010 7212 7630 7272
rect 9298 6848 10288 6900
rect 16942 6618 17798 6664
rect 14866 6418 15088 6472
rect 15696 6418 16176 6466
rect 11904 6300 13376 6348
rect 122 4756 166 5526
rect 14874 4574 15064 4654
rect 15812 4570 16102 4654
rect 17182 4268 17562 4366
rect 9404 3448 10264 3494
rect 12194 3436 13062 3498
rect 3256 2836 5312 2884
rect 6378 2848 8430 2896
rect 222 2726 960 2768
<< metal1 >>
rect -812 9296 19074 10100
rect -812 8898 -340 9296
rect 154 9142 1078 9296
rect 154 9102 246 9142
rect 982 9102 1078 9142
rect 154 9096 1078 9102
rect 1275 9038 1385 9039
rect 302 8988 1385 9038
rect -812 8392 302 8898
rect 1240 8820 1385 8988
rect 2003 8820 2121 8826
rect 1240 8812 2003 8820
rect 922 8702 2003 8812
rect 922 8582 1385 8702
rect 2003 8696 2121 8702
rect -812 7372 -340 8392
rect 1240 8308 1385 8582
rect 302 8258 1385 8308
rect 1275 7949 1385 8258
rect 1275 7839 1531 7949
rect 1422 7772 1530 7839
rect 1416 7664 1422 7772
rect 1530 7664 1536 7772
rect 2980 7590 3624 9296
rect 4634 8930 10692 9296
rect 4634 8882 4660 8930
rect 10668 8882 10692 8930
rect 4634 8876 10692 8882
rect 4075 8702 4081 8820
rect 4199 8774 10602 8820
rect 4199 8702 4404 8774
rect 11240 8746 11380 9296
rect 11733 8908 11871 9296
rect 11733 8792 11744 8908
rect 11860 8792 11871 8908
rect 11733 8781 11871 8792
rect 12044 8796 12580 9296
rect 4286 8292 4404 8702
rect 4662 8614 4672 8734
rect 4730 8614 4740 8734
rect 5978 8614 5988 8734
rect 6046 8614 6056 8734
rect 7292 8614 7302 8734
rect 7360 8614 7370 8734
rect 8610 8614 8620 8734
rect 8678 8614 8688 8734
rect 9924 8614 9934 8734
rect 9992 8614 10002 8734
rect 12044 8746 12072 8796
rect 12546 8746 12580 8796
rect 13754 8822 17860 9296
rect 13754 8774 13786 8822
rect 17822 8774 17860 8822
rect 13754 8768 17860 8774
rect 12044 8736 12580 8746
rect 13345 8712 13543 8713
rect 12140 8634 12836 8690
rect 11240 8600 11380 8606
rect 12078 8496 12088 8598
rect 12146 8496 12156 8598
rect 12334 8496 12344 8598
rect 12402 8496 12412 8598
rect 5320 8334 5330 8454
rect 5388 8334 5398 8454
rect 6634 8334 6644 8454
rect 6702 8334 6712 8454
rect 7952 8334 7962 8454
rect 8020 8334 8030 8454
rect 9268 8334 9278 8454
rect 9336 8334 9346 8454
rect 10584 8334 10594 8454
rect 10652 8334 10662 8454
rect 4286 8246 10602 8292
rect 12206 8266 12216 8368
rect 12274 8266 12284 8368
rect 12462 8266 12472 8368
rect 12530 8266 12540 8368
rect 12780 8238 12836 8634
rect 13345 8660 17756 8712
rect 12780 8228 13050 8238
rect 12140 8182 13050 8228
rect 13106 8182 13112 8238
rect 13345 8184 13554 8660
rect 18161 8632 18324 9296
rect 14444 8510 14454 8624
rect 14518 8510 14528 8624
rect 15760 8512 15770 8626
rect 15834 8512 15844 8626
rect 17076 8512 17086 8626
rect 17150 8512 17160 8626
rect 18161 8504 18178 8632
rect 18306 8504 18324 8632
rect 18161 8487 18324 8504
rect 13786 8226 13796 8340
rect 13860 8226 13870 8340
rect 15100 8226 15110 8340
rect 15174 8226 15184 8340
rect 16418 8226 16428 8340
rect 16492 8226 16502 8340
rect 17736 8226 17746 8340
rect 17810 8226 17820 8340
rect 12140 8172 12836 8182
rect 13345 8132 17756 8184
rect 12391 7959 12589 7965
rect 13345 7959 13543 8132
rect 12589 7761 13543 7959
rect 12391 7755 12589 7761
rect 7490 7590 9512 7594
rect -812 7364 180 7372
rect 1592 7368 1654 7369
rect -812 6584 126 7364
rect 166 6584 180 7364
rect 280 7306 1654 7368
rect 352 7170 362 7266
rect 418 7170 428 7266
rect 610 7170 620 7266
rect 676 7170 686 7266
rect 864 7170 874 7266
rect 930 7170 940 7266
rect 1120 7170 1130 7266
rect 1186 7170 1196 7266
rect 1414 6796 1530 6802
rect 1592 6796 1654 7306
rect 2979 7362 9512 7590
rect 2979 7272 7642 7362
rect 3984 7212 4010 7272
rect 7630 7212 7642 7272
rect 3984 7198 7642 7212
rect 7942 7168 8154 7170
rect 4052 7104 8154 7168
rect 3988 6964 3998 7070
rect 4056 6964 4066 7070
rect 4384 6964 4394 7070
rect 4452 6964 4462 7070
rect 4780 6964 4790 7070
rect 4848 6964 4858 7070
rect 5174 6964 5184 7070
rect 5242 6964 5252 7070
rect 5570 6964 5580 7070
rect 5638 6964 5648 7070
rect 5968 6964 5978 7070
rect 6036 6964 6046 7070
rect 6364 6964 6374 7070
rect 6432 6964 6442 7070
rect 6758 6964 6768 7070
rect 6826 6964 6836 7070
rect 7156 6964 7166 7070
rect 7224 6964 7234 7070
rect 7552 6964 7562 7070
rect 7620 6964 7630 7070
rect 238 6690 248 6786
rect 304 6690 314 6786
rect 482 6686 492 6782
rect 548 6686 558 6782
rect 736 6686 746 6782
rect 802 6686 812 6782
rect 994 6686 1004 6782
rect 1060 6686 1070 6782
rect 1530 6680 1654 6796
rect 4186 6772 4196 6878
rect 4254 6772 4264 6878
rect 4580 6772 4590 6878
rect 4648 6772 4658 6878
rect 4976 6772 4986 6878
rect 5044 6772 5054 6878
rect 5374 6772 5384 6878
rect 5442 6772 5452 6878
rect 5770 6772 5780 6878
rect 5838 6772 5848 6878
rect 6164 6772 6174 6878
rect 6232 6772 6242 6878
rect 6560 6772 6570 6878
rect 6628 6772 6638 6878
rect 6956 6772 6966 6878
rect 7024 6772 7034 6878
rect 7352 6772 7362 6878
rect 7420 6772 7430 6878
rect 7942 6726 8154 7104
rect 9280 7132 9512 7362
rect 13682 7270 17443 7474
rect 9280 6900 10312 7132
rect 9280 6848 9298 6900
rect 10288 6848 10312 6900
rect 9280 6842 10312 6848
rect 1414 6664 1654 6680
rect 1414 6636 1658 6664
rect 4056 6662 8154 6726
rect -812 6570 180 6584
rect 280 6574 1658 6636
rect -354 6568 180 6570
rect -854 5926 677 6239
rect 990 5926 996 6239
rect -326 5582 172 5584
rect -782 5526 172 5582
rect 1538 5538 1658 6574
rect 7942 5790 8154 6662
rect 8930 6736 10228 6790
rect 13682 6768 13886 7270
rect 18617 7026 18979 9296
rect 8930 6312 9064 6736
rect 11976 6718 13886 6768
rect 14836 6901 18979 7026
rect 14836 6853 17998 6901
rect 14836 6723 15357 6853
rect 15487 6796 17998 6853
rect 15487 6723 16204 6796
rect 14836 6720 16204 6723
rect 9304 6570 9314 6702
rect 9374 6570 9384 6702
rect 9560 6570 9570 6702
rect 9630 6570 9640 6702
rect 9816 6570 9826 6702
rect 9886 6570 9896 6702
rect 10072 6570 10082 6702
rect 10142 6570 10152 6702
rect 11910 6608 11920 6688
rect 11980 6608 11990 6688
rect 12826 6610 12836 6690
rect 12896 6610 12906 6690
rect 13544 6608 13886 6718
rect 14439 6703 16204 6720
rect 12368 6486 12378 6566
rect 12438 6486 12448 6566
rect 13284 6486 13294 6566
rect 13354 6486 13364 6566
rect 13544 6458 13662 6608
rect 14439 6557 14455 6703
rect 14601 6642 16204 6703
rect 14601 6557 15118 6642
rect 14439 6541 15118 6557
rect 11976 6408 13662 6458
rect 14836 6472 15118 6541
rect 14836 6418 14866 6472
rect 15088 6418 15118 6472
rect 14836 6406 15118 6418
rect 15666 6466 16204 6642
rect 16924 6747 17998 6796
rect 18152 6747 18979 6901
rect 16924 6664 18979 6747
rect 16924 6618 16942 6664
rect 17798 6618 17828 6664
rect 16924 6610 17828 6618
rect 15666 6418 15696 6466
rect 16176 6418 16204 6466
rect 15666 6404 16204 6418
rect 16568 6504 17736 6560
rect 8645 6178 8651 6312
rect 8785 6232 9064 6312
rect 9432 6272 9442 6404
rect 9502 6272 9512 6404
rect 9690 6272 9700 6404
rect 9760 6272 9770 6404
rect 9944 6270 9954 6402
rect 10014 6270 10024 6402
rect 10200 6272 10210 6404
rect 10270 6272 10280 6404
rect 15424 6362 15512 6364
rect 11876 6348 13410 6354
rect 11876 6300 11904 6348
rect 13376 6300 13410 6348
rect 14616 6304 15024 6362
rect 15424 6306 16102 6362
rect 8785 6178 10228 6232
rect 11876 6120 13986 6300
rect 7942 5789 8160 5790
rect 7942 5594 8173 5789
rect 13806 5737 13986 6120
rect 14312 6032 14448 6038
rect 14616 6032 14700 6304
rect 14876 6146 14886 6270
rect 14942 6146 14952 6270
rect 14448 5896 14700 6032
rect 14312 5890 14448 5896
rect 14616 5830 14700 5896
rect 15004 5872 15014 5996
rect 15070 5872 15080 5996
rect 15424 5830 15512 6306
rect 15702 6156 15712 6268
rect 15772 6156 15782 6268
rect 15958 6156 15968 6268
rect 16028 6156 16038 6268
rect 15832 5872 15842 5984
rect 15902 5872 15912 5984
rect 16088 5872 16098 5984
rect 16158 5872 16168 5984
rect 16568 5853 16702 6504
rect 16948 6348 16958 6468
rect 17018 6348 17028 6468
rect 17202 6348 17212 6468
rect 17272 6348 17282 6468
rect 17460 6348 17470 6468
rect 17530 6348 17540 6468
rect 17714 6348 17724 6468
rect 17784 6348 17794 6468
rect 17076 5876 17086 5996
rect 17146 5876 17156 5996
rect 17330 5876 17340 5996
rect 17400 5876 17410 5996
rect 17586 5876 17596 5996
rect 17656 5876 17666 5996
rect 14616 5829 15024 5830
rect 14614 5772 15024 5829
rect 15424 5828 15516 5830
rect 16564 5828 16706 5853
rect 15424 5772 16102 5828
rect 16564 5772 17736 5828
rect -782 4756 122 5526
rect 166 4756 172 5526
rect 366 5468 1658 5538
rect 4044 5530 8173 5594
rect 228 5342 238 5440
rect 296 5342 306 5440
rect 416 5342 426 5440
rect 484 5342 494 5440
rect 608 5342 618 5440
rect 676 5342 686 5440
rect 800 5342 810 5440
rect 868 5342 878 5440
rect 1538 5293 1658 5468
rect 3988 5406 3998 5488
rect 4056 5406 4066 5488
rect 4384 5406 4394 5488
rect 4452 5406 4462 5488
rect 4780 5406 4790 5488
rect 4848 5406 4858 5488
rect 5176 5406 5186 5488
rect 5244 5406 5254 5488
rect 5572 5406 5582 5488
rect 5640 5406 5650 5488
rect 5968 5406 5978 5488
rect 6036 5406 6046 5488
rect 6364 5406 6374 5488
rect 6432 5406 6442 5488
rect 6760 5406 6770 5488
rect 6828 5406 6838 5488
rect 7156 5406 7166 5488
rect 7224 5406 7234 5488
rect 7552 5406 7562 5488
rect 7620 5406 7630 5488
rect 1158 5179 1164 5293
rect 1278 5179 1658 5293
rect 4186 5210 4196 5292
rect 4254 5210 4264 5292
rect 4582 5210 4592 5292
rect 4650 5210 4660 5292
rect 4978 5210 4988 5292
rect 5046 5210 5056 5292
rect 5372 5210 5382 5292
rect 5440 5210 5450 5292
rect 5768 5210 5778 5292
rect 5836 5210 5846 5292
rect 6166 5210 6176 5292
rect 6234 5210 6244 5292
rect 6560 5210 6570 5292
rect 6628 5210 6638 5292
rect 6958 5210 6968 5292
rect 7026 5210 7036 5292
rect 7354 5210 7364 5292
rect 7422 5210 7432 5292
rect 320 4854 330 4952
rect 388 4854 398 4952
rect 512 4854 522 4952
rect 580 4854 590 4952
rect 704 4854 714 4952
rect 772 4854 782 4952
rect 896 4854 906 4952
rect 964 4854 974 4952
rect 1538 4808 1658 5179
rect 7942 5162 8173 5530
rect 4044 5098 8173 5162
rect 7942 5094 8173 5098
rect 8035 5001 8173 5094
rect 11084 5596 11392 5602
rect 8035 4863 8377 5001
rect 8515 4863 8521 5001
rect -782 4718 172 4756
rect 276 4738 1658 4808
rect 1538 4736 1658 4738
rect -782 3502 -310 4718
rect 1176 4386 1288 4392
rect 1288 4382 1650 4386
rect 1288 4274 1666 4382
rect 1176 4268 1288 4274
rect 1530 3922 1666 4274
rect 2168 4334 6178 4522
rect 10472 4341 10478 4487
rect 10624 4341 10630 4487
rect 2168 3922 2356 4334
rect 5990 3942 6178 4334
rect 2570 3922 5284 3924
rect 1530 3856 5284 3922
rect 5988 3866 8382 3942
rect 10478 3912 10624 4341
rect 1530 3736 2858 3856
rect 1530 3598 1666 3736
rect 290 3538 1666 3598
rect -782 2916 284 3502
rect 894 3220 978 3502
rect 894 3219 1144 3220
rect 1530 3219 1666 3538
rect 894 3053 1666 3219
rect 894 3052 1144 3053
rect 894 2922 978 3052
rect -782 2486 -310 2916
rect 1530 2878 1666 3053
rect 2570 2996 2858 3736
rect 3256 3684 3266 3810
rect 3330 3684 3340 3810
rect 4572 3684 4582 3810
rect 4646 3684 4656 3810
rect 5568 3178 5718 3184
rect 3910 3038 3920 3164
rect 3984 3038 3994 3164
rect 5232 3038 5242 3164
rect 5306 3038 5316 3164
rect 2570 2946 5244 2996
rect 292 2830 1666 2878
rect 3244 2884 5332 2890
rect 3244 2836 3256 2884
rect 5312 2836 5332 2884
rect 170 2768 1018 2774
rect 170 2726 222 2768
rect 960 2726 1018 2768
rect 170 2486 1018 2726
rect 3244 2486 5332 2836
rect 5568 2486 5718 3028
rect 5990 3008 6178 3866
rect 9462 3864 10632 3912
rect 10460 3844 10632 3864
rect 6372 3684 6382 3826
rect 6456 3684 6466 3826
rect 7686 3684 7696 3826
rect 7770 3684 7780 3826
rect 9408 3754 9418 3836
rect 9474 3754 9484 3836
rect 9926 3754 9936 3836
rect 9992 3754 10002 3836
rect 10460 3766 10491 3844
rect 10569 3766 10632 3844
rect 9130 3644 9136 3716
rect 9208 3644 9214 3716
rect 9136 3388 9208 3644
rect 9668 3636 9678 3718
rect 9734 3636 9744 3718
rect 10182 3634 10192 3716
rect 10248 3634 10258 3716
rect 10460 3604 10632 3766
rect 11084 3662 11392 5288
rect 11896 4809 11998 4815
rect 11896 3922 11998 4707
rect 11896 3868 12994 3922
rect 9462 3556 10632 3604
rect 11896 3610 11998 3868
rect 12460 3766 12470 3840
rect 12526 3766 12536 3840
rect 12976 3766 12986 3840
rect 13042 3766 13052 3840
rect 12202 3640 12212 3714
rect 12268 3640 12278 3714
rect 12718 3638 12728 3712
rect 12784 3638 12794 3712
rect 11896 3562 12994 3610
rect 9386 3494 10288 3500
rect 9386 3448 9404 3494
rect 10264 3448 10288 3494
rect 9386 3388 10288 3448
rect 9136 3316 10288 3388
rect 12158 3498 13098 3504
rect 12158 3436 12194 3498
rect 13062 3436 13098 3498
rect 12158 3317 13098 3436
rect 8754 3200 8914 3206
rect 7030 3048 7040 3190
rect 7114 3048 7124 3190
rect 8344 3048 8354 3190
rect 8428 3048 8438 3190
rect 5990 2958 8358 3008
rect 6334 2896 8454 2902
rect 6334 2848 6378 2896
rect 8430 2848 8454 2896
rect 6334 2486 8454 2848
rect 8754 2486 8914 3040
rect 9386 2486 10288 3316
rect 11713 3171 11719 3317
rect 11865 3171 13098 3317
rect 12158 2486 13098 3171
rect 13755 2486 14037 5737
rect 14614 5082 14700 5772
rect 15424 5513 15516 5772
rect 16564 5536 16706 5772
rect 15189 5497 15516 5513
rect 15189 5391 15204 5497
rect 15310 5391 15516 5497
rect 15189 5376 15516 5391
rect 15424 5180 15516 5376
rect 16264 5513 16706 5536
rect 16264 5383 16286 5513
rect 16416 5383 16706 5513
rect 16264 5361 16706 5383
rect 16564 5190 16706 5361
rect 18168 5443 18898 5488
rect 18168 5317 18213 5443
rect 18339 5317 18898 5443
rect 18168 5272 18898 5317
rect 15424 5122 16044 5180
rect 16564 5136 17408 5190
rect 14614 5024 15014 5082
rect 14614 4762 14700 5024
rect 14978 4912 14988 4994
rect 15042 4912 15052 4994
rect 14884 4794 14894 4876
rect 14948 4794 14958 4876
rect 15424 4766 15516 5122
rect 15822 5000 15832 5086
rect 15892 5000 15902 5086
rect 16012 5000 16022 5086
rect 16082 5000 16092 5086
rect 15918 4804 15928 4890
rect 15988 4804 15998 4890
rect 16564 4860 16706 5136
rect 17280 4994 17290 5096
rect 17356 4994 17366 5096
rect 17472 4994 17482 5096
rect 17548 4994 17558 5096
rect 14614 4756 15014 4762
rect 15424 4756 15948 4766
rect 14616 4704 15014 4756
rect 15426 4710 15948 4756
rect 14848 4654 15094 4666
rect 14848 4574 14874 4654
rect 15064 4574 15094 4654
rect 14848 4521 15094 4574
rect 14462 4503 15094 4521
rect 14462 4401 14479 4503
rect 14581 4492 15094 4503
rect 15784 4654 16126 4662
rect 15784 4570 15812 4654
rect 16102 4570 16126 4654
rect 15784 4492 16126 4570
rect 14581 4401 16126 4492
rect 14462 4384 16126 4401
rect 14848 4366 16126 4384
rect 16428 4649 16737 4860
rect 16428 4423 16469 4649
rect 16695 4476 16737 4649
rect 17184 4518 17194 4620
rect 17260 4518 17270 4620
rect 17376 4520 17386 4622
rect 17452 4520 17462 4622
rect 16695 4423 17504 4476
rect 16428 4422 17504 4423
rect 16428 4382 16737 4422
rect 14848 4262 15572 4366
rect 15676 4262 16126 4366
rect 14848 4178 16126 4262
rect 17152 4366 17590 4374
rect 17152 4268 17182 4366
rect 17562 4268 17590 4366
rect 17152 4191 18914 4268
rect 17152 4178 17830 4191
rect 14846 4065 17830 4178
rect 17956 4065 18914 4191
rect 14846 3936 18914 4065
rect 18582 2486 18914 3936
rect -784 1682 19074 2486
<< via1 >>
rect 2003 8702 2121 8820
rect 1422 7664 1530 7772
rect 4081 8702 4199 8820
rect 11744 8792 11860 8908
rect 4672 8614 4730 8734
rect 5988 8614 6046 8734
rect 7302 8614 7360 8734
rect 8620 8614 8678 8734
rect 9934 8614 9992 8734
rect 11240 8606 11380 8746
rect 12088 8496 12146 8598
rect 12344 8496 12402 8598
rect 5330 8334 5388 8454
rect 6644 8334 6702 8454
rect 7962 8334 8020 8454
rect 9278 8334 9336 8454
rect 10594 8334 10652 8454
rect 12216 8266 12274 8368
rect 12472 8266 12530 8368
rect 13050 8182 13106 8238
rect 14454 8510 14518 8624
rect 15770 8512 15834 8626
rect 17086 8512 17150 8626
rect 18178 8504 18306 8632
rect 13796 8226 13860 8340
rect 15110 8226 15174 8340
rect 16428 8226 16492 8340
rect 17746 8226 17810 8340
rect 12391 7761 12589 7959
rect 362 7170 418 7266
rect 620 7170 676 7266
rect 874 7170 930 7266
rect 1130 7170 1186 7266
rect 3998 6964 4056 7070
rect 4394 6964 4452 7070
rect 4790 6964 4848 7070
rect 5184 6964 5242 7070
rect 5580 6964 5638 7070
rect 5978 6964 6036 7070
rect 6374 6964 6432 7070
rect 6768 6964 6826 7070
rect 7166 6964 7224 7070
rect 7562 6964 7620 7070
rect 248 6690 304 6786
rect 492 6686 548 6782
rect 746 6686 802 6782
rect 1004 6686 1060 6782
rect 1414 6680 1530 6796
rect 4196 6772 4254 6878
rect 4590 6772 4648 6878
rect 4986 6772 5044 6878
rect 5384 6772 5442 6878
rect 5780 6772 5838 6878
rect 6174 6772 6232 6878
rect 6570 6772 6628 6878
rect 6966 6772 7024 6878
rect 7362 6772 7420 6878
rect 677 5926 990 6239
rect 15357 6723 15487 6853
rect 9314 6570 9374 6702
rect 9570 6570 9630 6702
rect 9826 6570 9886 6702
rect 10082 6570 10142 6702
rect 11920 6608 11980 6688
rect 12836 6610 12896 6690
rect 12378 6486 12438 6566
rect 13294 6486 13354 6566
rect 14455 6557 14601 6703
rect 17998 6747 18152 6901
rect 8651 6178 8785 6312
rect 9442 6272 9502 6404
rect 9700 6272 9760 6404
rect 9954 6270 10014 6402
rect 10210 6272 10270 6404
rect 14886 6146 14942 6270
rect 14312 5896 14448 6032
rect 15014 5872 15070 5996
rect 15712 6156 15772 6268
rect 15968 6156 16028 6268
rect 15842 5872 15902 5984
rect 16098 5872 16158 5984
rect 16958 6348 17018 6468
rect 17212 6348 17272 6468
rect 17470 6348 17530 6468
rect 17724 6348 17784 6468
rect 17086 5876 17146 5996
rect 17340 5876 17400 5996
rect 17596 5876 17656 5996
rect 238 5342 296 5440
rect 426 5342 484 5440
rect 618 5342 676 5440
rect 810 5342 868 5440
rect 3998 5406 4056 5488
rect 4394 5406 4452 5488
rect 4790 5406 4848 5488
rect 5186 5406 5244 5488
rect 5582 5406 5640 5488
rect 5978 5406 6036 5488
rect 6374 5406 6432 5488
rect 6770 5406 6828 5488
rect 7166 5406 7224 5488
rect 7562 5406 7620 5488
rect 1164 5179 1278 5293
rect 4196 5210 4254 5292
rect 4592 5210 4650 5292
rect 4988 5210 5046 5292
rect 5382 5210 5440 5292
rect 5778 5210 5836 5292
rect 6176 5210 6234 5292
rect 6570 5210 6628 5292
rect 6968 5210 7026 5292
rect 7364 5210 7422 5292
rect 330 4854 388 4952
rect 522 4854 580 4952
rect 714 4854 772 4952
rect 906 4854 964 4952
rect 11084 5288 11392 5596
rect 8377 4863 8515 5001
rect 1176 4274 1288 4386
rect 10478 4341 10624 4487
rect 3266 3684 3330 3810
rect 4582 3684 4646 3810
rect 3920 3038 3984 3164
rect 5242 3038 5306 3164
rect 5568 3028 5718 3178
rect 6382 3684 6456 3826
rect 7696 3684 7770 3826
rect 9418 3754 9474 3836
rect 9936 3754 9992 3836
rect 10491 3766 10569 3844
rect 9136 3644 9208 3716
rect 9678 3636 9734 3718
rect 10192 3634 10248 3716
rect 11896 4707 11998 4809
rect 12470 3766 12526 3840
rect 12986 3766 13042 3840
rect 12212 3640 12268 3714
rect 12728 3638 12784 3712
rect 7040 3048 7114 3190
rect 8354 3048 8428 3190
rect 8754 3040 8914 3200
rect 11719 3171 11865 3317
rect 15204 5391 15310 5497
rect 16286 5383 16416 5513
rect 18213 5317 18339 5443
rect 14988 4912 15042 4994
rect 14894 4794 14948 4876
rect 15832 5000 15892 5086
rect 16022 5000 16082 5086
rect 15928 4804 15988 4890
rect 17290 4994 17356 5096
rect 17482 4994 17548 5096
rect 14479 4401 14581 4503
rect 16469 4423 16695 4649
rect 17194 4518 17260 4620
rect 17386 4520 17452 4622
rect 15572 4262 15676 4366
rect 17830 4065 17956 4191
<< metal2 >>
rect 11744 8908 11860 8914
rect 4081 8820 4199 8826
rect 1997 8702 2003 8820
rect 2121 8702 4081 8820
rect 3873 7959 3991 8702
rect 4081 8696 4199 8702
rect 4660 8734 11240 8746
rect 4660 8614 4672 8734
rect 4730 8614 5988 8734
rect 6046 8614 7302 8734
rect 7360 8614 8620 8734
rect 8678 8614 9934 8734
rect 9992 8614 11240 8734
rect 4660 8606 11240 8614
rect 11380 8606 11386 8746
rect 11744 8608 11860 8792
rect 14454 8632 14518 8634
rect 15770 8632 15834 8636
rect 17086 8632 17150 8636
rect 18178 8632 18306 8638
rect 14436 8626 18178 8632
rect 14436 8624 15770 8626
rect 4672 8604 4730 8606
rect 5988 8604 6046 8606
rect 7302 8604 7360 8606
rect 8620 8604 8678 8606
rect 9934 8604 9992 8606
rect 11744 8598 12410 8608
rect 11744 8496 12088 8598
rect 12146 8496 12344 8598
rect 12402 8496 12410 8598
rect 14436 8510 14454 8624
rect 14518 8512 15770 8624
rect 15834 8512 17086 8626
rect 17150 8512 18178 8626
rect 14518 8510 18178 8512
rect 14436 8504 18178 8510
rect 14454 8500 14518 8504
rect 15770 8502 15834 8504
rect 17086 8502 17150 8504
rect 18178 8498 18306 8504
rect 11744 8492 12410 8496
rect 12088 8486 12146 8492
rect 12344 8486 12402 8492
rect 5310 8454 11380 8466
rect 5310 8334 5330 8454
rect 5388 8334 6644 8454
rect 6702 8334 7962 8454
rect 8020 8334 9278 8454
rect 9336 8334 10594 8454
rect 10652 8334 11380 8454
rect 12216 8376 12274 8378
rect 12472 8376 12530 8378
rect 5310 8326 11380 8334
rect 5330 8324 5388 8326
rect 6644 8324 6702 8326
rect 7962 8324 8020 8326
rect 9278 8324 9336 8326
rect 10594 8324 10652 8326
rect 1422 7772 1530 7778
rect 3833 7761 10121 7959
rect 10319 7761 10328 7959
rect 362 7272 418 7276
rect 620 7272 676 7276
rect 874 7272 930 7276
rect 1130 7272 1186 7276
rect 1422 7272 1530 7664
rect 350 7266 1530 7272
rect 350 7170 362 7266
rect 418 7170 620 7266
rect 676 7170 874 7266
rect 930 7170 1130 7266
rect 1186 7170 1530 7266
rect 350 7164 1530 7170
rect 8957 7455 10825 7457
rect 11012 7455 11380 8326
rect 8957 7355 11380 7455
rect 362 7160 418 7164
rect 620 7160 676 7164
rect 874 7160 930 7164
rect 1130 7160 1186 7164
rect 2519 7078 3262 7168
rect 3998 7078 4056 7080
rect 4394 7078 4452 7080
rect 4790 7078 4848 7080
rect 5184 7078 5242 7080
rect 5580 7078 5638 7080
rect 5978 7078 6036 7080
rect 6374 7078 6432 7080
rect 6768 7078 6826 7080
rect 7166 7078 7224 7080
rect 7562 7078 7620 7080
rect 2519 7070 7627 7078
rect 2519 6964 3998 7070
rect 4056 6964 4394 7070
rect 4452 6964 4790 7070
rect 4848 6964 5184 7070
rect 5242 6964 5580 7070
rect 5638 6964 5978 7070
rect 6036 6964 6374 7070
rect 6432 6964 6768 7070
rect 6826 6964 7166 7070
rect 7224 6964 7562 7070
rect 7620 6964 7627 7070
rect 2519 6944 7627 6964
rect 2519 6855 3262 6944
rect 4196 6882 4254 6888
rect 4590 6882 4648 6888
rect 4986 6882 5044 6888
rect 5384 6882 5442 6888
rect 5780 6882 5838 6888
rect 6174 6882 6232 6888
rect 6570 6882 6628 6888
rect 6966 6882 7024 6888
rect 7362 6882 7420 6888
rect 3430 6878 7444 6882
rect 246 6786 1414 6796
rect 246 6690 248 6786
rect 304 6782 1414 6786
rect 304 6690 492 6782
rect 246 6686 492 6690
rect 548 6686 746 6782
rect 802 6686 1004 6782
rect 1060 6686 1414 6782
rect 246 6680 1414 6686
rect 1530 6680 1536 6796
rect 492 6676 548 6680
rect 746 6676 802 6680
rect 1004 6676 1060 6680
rect 677 6239 990 6245
rect 2519 6239 2832 6855
rect 3430 6772 4196 6878
rect 4254 6772 4590 6878
rect 4648 6772 4986 6878
rect 5044 6772 5384 6878
rect 5442 6772 5780 6878
rect 5838 6772 6174 6878
rect 6232 6772 6570 6878
rect 6628 6772 6966 6878
rect 7024 6772 7362 6878
rect 7420 6772 7444 6878
rect 3430 6764 7444 6772
rect 990 5926 2832 6239
rect 3435 6312 3577 6764
rect 4196 6762 4254 6764
rect 4590 6762 4648 6764
rect 4986 6762 5044 6764
rect 5384 6762 5442 6764
rect 5780 6762 5838 6764
rect 6174 6762 6232 6764
rect 6570 6762 6628 6764
rect 6966 6762 7024 6764
rect 7362 6762 7420 6764
rect 8957 6712 9059 7355
rect 10711 7353 11380 7355
rect 11012 7352 11380 7353
rect 11648 8368 12534 8376
rect 11648 8266 12216 8368
rect 12274 8266 12472 8368
rect 12530 8266 12534 8368
rect 13784 8340 18170 8350
rect 11648 8254 12534 8266
rect 8957 6702 10172 6712
rect 8957 6570 9314 6702
rect 9374 6570 9570 6702
rect 9630 6570 9826 6702
rect 9886 6570 10082 6702
rect 10142 6570 10172 6702
rect 11090 6570 11379 7352
rect 11648 6698 11738 8254
rect 13016 8238 13141 8273
rect 13016 8182 13050 8238
rect 13106 8182 13141 8238
rect 13784 8226 13796 8340
rect 13860 8226 15110 8340
rect 15174 8226 16428 8340
rect 16492 8226 17746 8340
rect 17810 8226 18170 8340
rect 13784 8212 18170 8226
rect 12102 7959 12290 7963
rect 12097 7954 12391 7959
rect 12097 7766 12102 7954
rect 12290 7766 12391 7954
rect 12097 7761 12391 7766
rect 12589 7761 12595 7959
rect 12102 7757 12290 7761
rect 12104 7245 12113 7471
rect 12339 7421 12881 7471
rect 13016 7421 13141 8182
rect 18032 7921 18170 8212
rect 14189 7783 18170 7921
rect 14189 7522 14327 7783
rect 12339 7296 13141 7421
rect 14186 7413 14327 7522
rect 12339 7245 12881 7296
rect 14186 7002 14322 7413
rect 14068 6866 14322 7002
rect 17998 6901 18152 6907
rect 12836 6698 12896 6700
rect 11648 6690 12916 6698
rect 11648 6688 12836 6690
rect 11648 6608 11920 6688
rect 11980 6610 12836 6688
rect 12896 6610 12916 6690
rect 11980 6608 12916 6610
rect 11920 6598 11980 6608
rect 12836 6600 12896 6608
rect 8957 6558 10172 6570
rect 11084 6566 11392 6570
rect 12378 6566 12438 6576
rect 13294 6566 13354 6576
rect 8651 6312 8785 6318
rect 3435 6178 8651 6312
rect 677 5920 990 5926
rect 3435 5517 3577 6178
rect 8651 6172 8785 6178
rect 238 5440 1278 5450
rect 296 5342 426 5440
rect 484 5342 618 5440
rect 676 5342 810 5440
rect 868 5342 1278 5440
rect 238 5336 1278 5342
rect 238 5332 296 5336
rect 426 5332 484 5336
rect 618 5332 676 5336
rect 810 5332 868 5336
rect 1164 5293 1278 5336
rect 1164 5173 1278 5179
rect 2818 5375 3577 5517
rect 8957 5500 9059 6558
rect 11084 6486 12378 6566
rect 12438 6486 13294 6566
rect 13354 6486 13362 6566
rect 11084 6474 13362 6486
rect 9432 6404 10624 6420
rect 9432 6274 9442 6404
rect 9502 6274 9700 6404
rect 9442 6262 9502 6272
rect 9760 6402 10210 6404
rect 9760 6274 9954 6402
rect 9700 6262 9760 6272
rect 10014 6274 10210 6402
rect 9954 6260 10014 6270
rect 10270 6274 10624 6404
rect 10210 6262 10270 6272
rect 3988 5488 9059 5500
rect 3988 5406 3998 5488
rect 4056 5406 4394 5488
rect 4452 5406 4790 5488
rect 4848 5406 5186 5488
rect 5244 5406 5582 5488
rect 5640 5406 5978 5488
rect 6036 5406 6374 5488
rect 6432 5406 6770 5488
rect 6828 5406 7166 5488
rect 7224 5406 7562 5488
rect 7620 5406 9059 5488
rect 3988 5398 9059 5406
rect 3998 5396 4056 5398
rect 4394 5396 4452 5398
rect 4790 5396 4848 5398
rect 5186 5396 5244 5398
rect 5582 5396 5640 5398
rect 5978 5396 6036 5398
rect 6374 5396 6432 5398
rect 6770 5396 6828 5398
rect 7166 5396 7224 5398
rect 7562 5396 7620 5398
rect 330 4952 1288 4962
rect 388 4854 522 4952
rect 580 4854 714 4952
rect 772 4854 906 4952
rect 964 4854 1288 4952
rect 330 4850 1288 4854
rect 330 4844 388 4850
rect 522 4844 580 4850
rect 714 4844 772 4850
rect 906 4844 964 4850
rect 1176 4386 1288 4850
rect 1170 4274 1176 4386
rect 1288 4274 1294 4386
rect 2818 3816 2960 5375
rect 8344 5320 8556 5326
rect 8716 5320 8876 5334
rect 4156 5292 8876 5320
rect 4156 5210 4196 5292
rect 4254 5210 4592 5292
rect 4650 5210 4988 5292
rect 5046 5210 5382 5292
rect 5440 5210 5778 5292
rect 5836 5210 6176 5292
rect 6234 5210 6570 5292
rect 6628 5210 6968 5292
rect 7026 5210 7364 5292
rect 7422 5210 8876 5292
rect 4156 5188 8876 5210
rect 8377 5001 8515 5188
rect 8377 4857 8515 4863
rect 6382 3830 6456 3836
rect 7696 3830 7770 3836
rect 8716 3830 8876 5188
rect 10478 4839 10624 6274
rect 11084 5596 11392 6474
rect 14068 6032 14204 6866
rect 15357 6853 15487 6859
rect 14455 6703 14601 6709
rect 14455 6282 14601 6557
rect 14455 6270 14942 6282
rect 14455 6146 14886 6270
rect 15357 6278 15487 6723
rect 17998 6480 18152 6747
rect 16946 6468 18152 6480
rect 16946 6348 16958 6468
rect 17018 6348 17212 6468
rect 17272 6348 17470 6468
rect 17530 6348 17724 6468
rect 17784 6348 18152 6468
rect 16946 6326 18152 6348
rect 15357 6268 16032 6278
rect 15357 6156 15712 6268
rect 15772 6156 15968 6268
rect 16028 6156 16032 6268
rect 15357 6148 16032 6156
rect 15712 6146 15772 6148
rect 15968 6146 16028 6148
rect 14455 6136 14942 6146
rect 13398 6030 13656 6032
rect 14068 6030 14312 6032
rect 13398 5896 14312 6030
rect 14448 5896 14454 6032
rect 15012 5996 15310 6006
rect 13398 5894 14204 5896
rect 11078 5288 11084 5596
rect 11392 5288 11398 5596
rect 10478 4809 12028 4839
rect 10478 4707 11896 4809
rect 11998 4707 12028 4809
rect 10478 4678 12028 4707
rect 10478 4487 10624 4678
rect 10478 4335 10624 4341
rect 13398 3850 13656 5894
rect 15012 5872 15014 5996
rect 15070 5872 15310 5996
rect 17084 5996 18154 6008
rect 15842 5992 15902 5994
rect 16098 5992 16158 5994
rect 15012 5860 15310 5872
rect 15834 5984 16416 5992
rect 15834 5872 15842 5984
rect 15902 5872 16098 5984
rect 16158 5872 16416 5984
rect 15834 5862 16416 5872
rect 17084 5876 17086 5996
rect 17146 5876 17340 5996
rect 17400 5876 17596 5996
rect 17656 5876 18154 5996
rect 17084 5866 18154 5876
rect 15204 5497 15310 5860
rect 16286 5513 16416 5862
rect 15204 5008 15310 5391
rect 16280 5383 16286 5513
rect 16416 5383 16422 5513
rect 18028 5443 18154 5866
rect 16286 5096 16416 5383
rect 18028 5317 18213 5443
rect 18339 5317 18345 5443
rect 18028 5106 18154 5317
rect 17288 5096 18154 5106
rect 14988 4994 15310 5008
rect 15828 5086 16420 5096
rect 15828 5000 15832 5086
rect 15892 5000 16022 5086
rect 16082 5000 16420 5086
rect 15828 4996 16420 5000
rect 15042 4912 15310 4994
rect 15832 4990 15892 4996
rect 16022 4990 16082 4996
rect 16286 4995 16416 4996
rect 17288 4994 17290 5096
rect 17356 4994 17482 5096
rect 17548 4994 18154 5096
rect 17288 4980 18154 4994
rect 14988 4902 15310 4912
rect 15928 4898 15988 4900
rect 15572 4890 15994 4898
rect 14479 4876 14948 4886
rect 14479 4794 14894 4876
rect 14479 4784 14948 4794
rect 15572 4804 15928 4890
rect 15988 4804 15994 4890
rect 15572 4794 15994 4804
rect 14479 4503 14581 4784
rect 14479 4395 14581 4401
rect 15572 4366 15676 4794
rect 15572 4256 15676 4262
rect 16469 4649 16695 4655
rect 17184 4622 17956 4632
rect 17184 4620 17386 4622
rect 17184 4518 17194 4620
rect 17260 4520 17386 4620
rect 17452 4520 17956 4622
rect 17260 4518 17956 4520
rect 17184 4506 17956 4518
rect 6360 3826 8876 3830
rect 3266 3816 3330 3820
rect 4582 3816 4646 3820
rect 2818 3810 4726 3816
rect 2818 3684 3266 3810
rect 3330 3684 4582 3810
rect 4646 3684 4726 3810
rect 2818 3674 4726 3684
rect 6360 3684 6382 3826
rect 6456 3684 7696 3826
rect 7770 3684 8876 3826
rect 9418 3844 9474 3846
rect 9936 3844 9992 3846
rect 9418 3836 10491 3844
rect 9474 3766 9936 3836
rect 9418 3744 9474 3754
rect 9992 3766 10491 3836
rect 10569 3766 10575 3844
rect 12464 3840 13656 3850
rect 12464 3766 12470 3840
rect 12526 3766 12986 3840
rect 13042 3836 13656 3840
rect 13042 3766 13651 3836
rect 12464 3760 13651 3766
rect 12470 3756 12526 3760
rect 12986 3756 13042 3760
rect 9936 3744 9992 3754
rect 6360 3670 8876 3684
rect 9136 3716 9208 3722
rect 9678 3718 9734 3728
rect 9208 3644 9678 3716
rect 9136 3638 9208 3644
rect 10192 3716 10248 3726
rect 12212 3722 12268 3724
rect 9734 3644 10192 3716
rect 9678 3626 9734 3636
rect 10248 3644 10250 3716
rect 11746 3714 12790 3722
rect 10192 3624 10248 3634
rect 11746 3640 12212 3714
rect 12268 3712 12790 3714
rect 12268 3640 12728 3712
rect 11746 3638 12728 3640
rect 12784 3638 12790 3712
rect 11746 3630 12790 3638
rect 11746 3459 11838 3630
rect 12728 3628 12784 3630
rect 16469 3512 16695 4423
rect 17830 4191 17956 4506
rect 17830 4059 17956 4065
rect 11719 3317 11865 3459
rect 7018 3190 8754 3200
rect 3906 3164 5568 3178
rect 3906 3038 3920 3164
rect 3984 3038 5242 3164
rect 5306 3038 5568 3164
rect 3906 3028 5568 3038
rect 5718 3028 5724 3178
rect 7018 3048 7040 3190
rect 7114 3048 8354 3190
rect 8428 3048 8754 3190
rect 7018 3040 8754 3048
rect 8914 3040 8920 3200
rect 16469 3296 16474 3512
rect 16690 3296 16695 3512
rect 16469 3291 16695 3296
rect 16474 3287 16690 3291
rect 11719 3165 11865 3171
rect 7040 3038 7114 3040
rect 8354 3038 8428 3040
<< via2 >>
rect 10121 7761 10319 7959
rect 12102 7766 12290 7954
rect 12113 7245 12339 7471
rect 16474 3296 16690 3512
<< metal3 >>
rect 10116 7959 10324 7964
rect 10116 7761 10121 7959
rect 10319 7954 12295 7959
rect 10319 7766 12102 7954
rect 12290 7766 12295 7954
rect 10319 7761 12295 7766
rect 10116 7756 10324 7761
rect 12108 7471 12344 7476
rect 11337 7245 12113 7471
rect 12339 7245 12344 7471
rect 11337 5967 11563 7245
rect 12108 7240 12344 7245
rect 11337 5741 12911 5967
rect 12685 4773 12911 5741
rect 12685 4547 14091 4773
rect 13865 3517 14091 4547
rect 13865 3512 16695 3517
rect 13865 3296 16474 3512
rect 16690 3296 16695 3512
rect 13865 3291 16695 3296
use sky130_fd_pr__nfet_01v8_lvt_BSZA4P  XM1
timestamp 1716907293
transform 1 0 12628 0 1 3740
box -554 -310 554 310
use sky130_fd_pr__nfet_01v8_lvt_BSZA4P  XM2
timestamp 1716907293
transform 1 0 9834 0 1 3734
box -554 -310 554 310
use sky130_fd_pr__pfet_01v8_lvt_366EDY  XM3
timestamp 1716907293
transform 1 0 9793 0 1 6485
box -615 -433 615 433
use sky130_fd_pr__pfet_01v8_lvt_ET6TZU  XM4
timestamp 1716907293
transform 1 0 5809 0 1 5349
box -1949 -369 1949 369
use sky130_fd_pr__pfet_01v8_lvt_ET6TZU  XM5
timestamp 1716907293
transform 1 0 5809 0 1 6915
box -1949 -369 1949 369
use sky130_fd_pr__pfet_01v8_lvt_CE5TV5  XM6
timestamp 1716907293
transform 1 0 7662 0 1 8533
box -3128 -419 3128 419
use sky130_fd_pr__pfet_01v8_lvt_QBWM73  XM7
timestamp 1716907293
transform 1 0 12309 0 1 8430
box -359 -386 359 386
use sky130_fd_pr__nfet_01v8_lvt_XWWVRJ  XM8
timestamp 1716907293
transform 1 0 12638 0 1 6588
box -854 -310 854 310
use sky130_fd_pr__pfet_01v8_lvt_CEZKS5  XM9
timestamp 1716907293
transform 1 0 15803 0 1 8423
box -2141 -419 2141 419
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XM10
timestamp 1716907293
transform 1 0 14969 0 1 4894
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_lvt_4QFWD3  XM11
timestamp 1716907293
transform 1 0 14979 0 1 6069
box -231 -419 231 419
use sky130_fd_pr__pfet_01v8_lvt_4QPJD3  XM12
timestamp 1716907293
transform 1 0 15935 0 1 6069
box -359 -419 359 419
use sky130_fd_pr__nfet_01v8_lvt_CW7PBK  XM13
timestamp 1716907293
transform 1 0 15957 0 1 4944
box -263 -360 263 360
use sky130_fd_pr__pfet_01v8_lvt_4QK4B3  XM14
timestamp 1716907293
transform 1 0 17371 0 1 6169
box -551 -519 551 519
use sky130_fd_pr__nfet_01v8_lvt_E5PS5K  XM15
timestamp 1716907293
transform 1 0 17371 0 1 4806
box -311 -510 311 510
use sky130_fd_pr__nfet_01v8_lvt_HEVHEL  XM16
timestamp 1716907293
transform 1 0 7404 0 1 3436
box -1154 -610 1154 610
use sky130_fd_pr__nfet_01v8_lvt_HEVHEL  XM17
timestamp 1716907293
transform 1 0 4284 0 1 3424
box -1154 -610 1154 610
use sky130_fd_pr__nfet_01v8_lvt_UJF2WX  XM18
timestamp 1716907293
transform 1 0 592 0 1 3208
box -496 -510 496 510
use sky130_fd_pr__pfet_01v8_lvt_CEYSV5  XM19
timestamp 1716907293
transform 1 0 614 0 1 8653
box -496 -519 496 519
use sky130_fd_pr__nfet_01v8_lvt_95PS5T  XM20
timestamp 1716907293
transform 1 0 599 0 1 5140
box -503 -510 503 510
use sky130_fd_pr__pfet_01v8_lvt_4QPHR2  XM21
timestamp 1716907293
transform 1 0 711 0 1 6975
box -615 -519 615 519
<< labels >>
flabel metal1 -704 1944 -504 2144 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 -798 5982 -598 6182 0 FreeSans 256 0 0 0 vref
port 2 nsew
flabel metal1 1530 3736 2638 3922 0 FreeSans 1600 0 0 0 i_n
flabel metal1 1538 4736 1658 6664 0 FreeSans 1600 0 0 0 dcon
flabel metal2 3435 5375 3577 6882 0 FreeSans 1600 0 0 0 vm
flabel metal2 8716 3670 8876 5334 0 FreeSans 1600 0 0 0 g1
flabel metal2 2121 8702 4081 8820 0 FreeSans 1600 0 0 0 vgb
flabel metal1 18694 5274 18894 5474 0 FreeSans 256 0 0 0 out
port 4 nsew
flabel metal1 11138 3716 11338 3916 0 FreeSans 256 0 0 0 in
port 5 nsew
flabel metal2 10478 4678 11896 4839 0 FreeSans 1600 0 0 0 g2
flabel metal2 14189 7783 18170 7921 0 FreeSans 1600 0 0 0 out1
flabel metal1 -686 9592 -486 9792 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 15424 4756 15516 5830 0 FreeSans 1600 0 0 0 out2
flabel metal1 16568 4422 16702 6560 0 FreeSans 1600 0 0 0 out3
flabel metal1 17235 7270 17435 7470 0 FreeSans 256 90 0 0 vgf
port 3 nsew
<< end >>

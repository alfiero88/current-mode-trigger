** sch_path: /home/ttuser/tt07-current-mode-trigger/xschem/CurrentTrigger.sch
.subckt CurrentTrigger vdd vss vref vgf out in
*.PININFO vdd:B vss:B in:I out:O vref:I vgf:I
XM1 out1 g2 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=3 m=1
XM2 g2 g2 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=3 m=1
XM3 g2 vm in vdd sky130_fd_pr__pfet_01v8_lvt L=0.35 W=15 nf=7 m=1
XM4 g1 g1 in vdd sky130_fd_pr__pfet_01v8_lvt L=0.7 W=27 nf=18 m=1
XM5 vm g1 vref vdd sky130_fd_pr__pfet_01v8_lvt L=0.7 W=27 nf=18 m=1
XM6 in vgb vdd vdd sky130_fd_pr__pfet_01v8_lvt L=3 W=18 nf=9 m=1
XM7 net1 out3 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.35 W=5 nf=5 m=1
XM9 out1 vgb vdd vdd sky130_fd_pr__pfet_01v8_lvt L=3 W=12 nf=6 m=1
XM10 out2 out1 vss vss sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 m=1
XM11 out2 out1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.35 W=2 nf=1 m=1
XM12 out3 out2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.35 W=6 nf=3 m=1
XM13 out3 out2 vss vss sky130_fd_pr__nfet_01v8_lvt L=0.15 W=3 nf=2 m=1
XM14 out out3 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.35 W=18 nf=6 m=1
XM15 out out3 vss vss sky130_fd_pr__nfet_01v8_lvt L=0.15 W=9 nf=3 m=1
XM16 g1 i_n vss vss sky130_fd_pr__nfet_01v8_lvt L=3 W=12 nf=3 m=1
XM17 vm i_n vss vss sky130_fd_pr__nfet_01v8_lvt L=3 W=12 nf=3 m=1
XM18 i_n i_n vss vss sky130_fd_pr__nfet_01v8_lvt L=3 W=3 nf=1 m=1
XM19 vgb vgb vdd vdd sky130_fd_pr__pfet_01v8_lvt L=3 W=3 nf=1 m=1
XM20 dcon dcon i_n vss sky130_fd_pr__nfet_01v8_lvt L=0.15 W=21 nf=7 m=1
XM21 dcon dcon vgb vdd sky130_fd_pr__pfet_01v8_lvt L=0.35 W=21 nf=7 m=1
XM8 net1 vgf in vss sky130_fd_pr__nfet_01v8_lvt L=2 W=3 nf=3 m=1
.ends
.end
